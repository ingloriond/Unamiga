LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;
PACKAGE rom_pack IS

  TYPE arr16 IS ARRAY(natural RANGE<>) OF unsigned(15 DOWNTO 0);
  TYPE arr8  IS ARRAY(natural RANGE<>) OF unsigned(7 DOWNTO 0);

  CONSTANT INIT_EXEC : arr16 := (
    x"0004",x"0112",x"0026",x"00AF",x"0270",x"0030",x"0270",x"0271",
    x"0272",x"0034",x"0273",x"0274",x"0275",x"00BD",x"02FD",x"0006",
    x"02BC",x"0100",x"0001",x"02A7",x"02B5",x"02B4",x"02B3",x"02B2",
    x"02B1",x"02B0",x"0038",x"02B0",x"02B7",x"02A9",x"0041",x"0288",
    x"0040",x"03B8",x"00FC",x"022C",x"0021",x"008F",x"02BE",x"02F1",
    x"0004",x"0118",x"0283",x"02B8",x"0026",x"0240",x"0100",x"02B8",
    x"0011",x"0240",x"0101",x"0001",x"02B8",x"0014",x"0050",x"0240",
    x"02F0",x"0004",x"0110",x"001D",x"0070",x"0004",x"0110",x"001D",
    x"0048",x"02B8",x"00FE",x"02BC",x"0102",x"0004",x"0114",x"0338",
    x"0004",x"0110",x"0060",x"035E",x"03FF",x"0147",x"0001",x"0115",
    x"000C",x"0116",x"00A0",x"0117",x"0008",x"0118",x"0060",x"0119",
    x"0008",x"0104",x"0008",x"0102",x"0084",x"0000",x"02A8",x"0248",
    x"02A9",x"0089",x"022C",x"0005",x"0002",x"0340",x"0102",x"0224",
    x"0003",x"0004",x"011C",x"0238",x"0004",x"0116",x"03B3",x"0004",
    x"0114",x"03FE",x"02B8",x"0090",x"0240",x"0102",x"0001",x"02B8",
    x"0006",x"0019",x"0240",x"035D",x"0004",x"0114",x"00F1",x"0004",
    x"0114",x"001C",x"0004",x"0110",x"00AB",x"000E",x"0245",x"0105",
    x"033C",x"000B",x"00BD",x"02FD",x"0004",x"0001",x"02A7",x"0002",
    x"0280",x"0102",x"0010",x"0223",x"0005",x"0281",x"0103",x"0241",
    x"0102",x"0020",x"0004",x"0114",x"027D",x"0004",x"0110",x"01FA",
    x"0004",x"0114",x"03D5",x"0004",x"0114",x"00F1",x"0004",x"0118",
    x"02AD",x"0220",x"001B",x"02AC",x"0275",x"037C",x"000C",x"020D",
    x"0007",x"02C4",x"02F0",x"033C",x"0014",x"0001",x"02A5",x"02B7",
    x"02C4",x"02F0",x"033C",x"0014",x"02A5",x"02B7",x"007D",x"0201",
    x"003F",x"0202",x"0013",x"007D",x"0201",x"003B",x"0202",x"0086",
    x"007D",x"0201",x"003C",x"0202",x"0051",x"02B9",x"0080",x"0241",
    x"002C",x"0009",x"0241",x"0102",x"0200",x"0028",x"0285",x"0021",
    x"01ED",x"02BC",x"0030",x"0265",x"0265",x"0265",x"02B8",x"000B",
    x"0240",x"0028",x"0240",x"002C",x"0268",x"037D",x"0008",x"022C",
    x"0004",x"0001",x"02B9",x"00A8",x"0036",x"02BB",x"0007",x"02BC",
    x"023D",x"0004",x"011A",x"0067",x"00A9",x"02BC",x"02C9",x"0004",
    x"0118",x"0067",x"02B8",x"0088",x"0240",x"0102",x"0240",x"0020",
    x"02B7",x"0241",x"0102",x"0004",x"011E",x"032F",x"02B7",x"0004",
    x"0110",x"00AB",x"000D",x"0245",x"0032",x"02A0",x"0078",x"0280",
    x"0021",x"0209",x"0002",x"0240",x"0021",x"02B9",x"0028",x"02B8",
    x"0005",x"0004",x"0114",x"0330",x"0241",x"0106",x"0281",x"0106",
    x"0241",x"002C",x"02B8",x"0003",x"0220",x"0029",x"0275",x"0281",
    x"0102",x"0041",x"0041",x"022B",x"006E",x"0011",x"020B",x"001E",
    x"0241",x"0102",x"0379",x"0003",x"020D",x"0018",x"0004",x"0110",
    x"0154",x"0280",x"0114",x"0080",x"0204",x"0006",x"03C0",x"0102",
    x"020C",x"000C",x"0240",x"0114",x"0240",x"0020",x"0004",x"0110",
    x"01C0",x"0004",x"0114",x"0014",x"0200",x"0002",x"0240",x"0020",
    x"02B5",x"0004",x"0318",x"02BD",x"0275",x"0049",x"00CF",x"0200",
    x"0052",x"0200",x"0006",x"01ED",x"02BC",x"031D",x"01DB",x"0200",
    x"0006",x"02BD",x"0004",x"02BC",x"033D",x"02BB",x"0004",x"02A0",
    x"0081",x"0065",x"0065",x"03B9",x"0380",x"0049",x"02A2",x"0092",
    x"02A2",x"0204",x"0004",x"0343",x"0104",x"0205",x"0003",x"02BA",
    x"00FF",x"000F",x"0042",x"03BA",x"00FF",x"01D1",x"0269",x"0081",
    x"0061",x"03B9",x"03E0",x"004D",x"02A2",x"0042",x"03BA",x"007F",
    x"01D1",x"02FD",x"0007",x"0269",x"0081",x"03B8",x"0007",x"03B9",
    x"0030",x"03F9",x"0008",x"0041",x"01C1",x"009A",x"02C2",x"02F0",
    x"03D1",x"02FD",x"0007",x"0269",x"02FD",x"0007",x"01C0",x"0268",
    x"02FC",x"0004",x"033D",x"0018",x"000B",x"0098",x"03B8",x"0003",
    x"022C",x"0042",x"02B7",x"02BC",x"0018",x"02BD",x"0107",x"02A0",
    x"0268",x"0040",x"0070",x"0034",x"0072",x"0070",x"0073",x"037D",
    x"010F",x"022C",x"000B",x"0042",x"026A",x"0043",x"026B",x"02B7",
    x"0275",x"0284",x"0112",x"0282",x"0111",x"007E",x"0004",x"0110",
    x"01D1",x"0284",x"0113",x"0282",x"0111",x"0062",x"007A",x"000A",
    x"000F",x"0275",x"0014",x"022B",x"00D4",x"01C9",x"0029",x"00E4",
    x"00E4",x"00E4",x"0285",x"02F0",x"00EA",x"033D",x"0014",x"0001",
    x"02EC",x"0295",x"0001",x"02FD",x"0000",x"0038",x"02A0",x"0268",
    x"02A0",x"0268",x"02A0",x"0268",x"02A0",x"0268",x"02A0",x"0268",
    x"02A0",x"0268",x"02A0",x"0268",x"02A0",x"0268",x"0011",x"0224",
    x"0012",x"02B7",x"0275",x"01C0",x"02B9",x"031D",x"02BA",x"0001",
    x"0200",x"001F",x"0240",x"011B",x"0241",x"031B",x"0242",x"011C",
    x"0004",x"0110",x"0226",x"002F",x"0012",x"0004",x"0110",x"0226",
    x"000B",x"0013",x"0004",x"0110",x"0226",x"00F9",x"0013",x"0282",
    x"011C",x"004A",x"0281",x"031B",x"02F9",x"0008",x"0280",x"011B",
    x"0008",x"0340",x"0104",x"0225",x"0022",x"02B7",x"0281",x"031B",
    x"0009",x"028C",x"00A4",x"0224",x"0015",x"0001",x"02AF",x"0275",
    x"0244",x"0319",x"02A1",x"03B9",x"0300",x"020C",x"0012",x"0280",
    x"011C",x"0380",x"0110",x"0204",x"000C",x"0274",x"0014",x"0001",
    x"03E1",x"0204",x"0005",x"0241",x"031C",x"0004",x"0114",x"00A1",
    x"02B4",x"02FC",x"0005",x"02A0",x"0078",x"0209",x"0012",x"0001",
    x"02A2",x"0281",x"011C",x"0381",x"010F",x"0204",x"0009",x"0242",
    x"031C",x"0270",x"0274",x"0004",x"0114",x"00A1",x"02B4",x"02B0",
    x"0080",x"0224",x"003D",x"0281",x"011B",x"02F9",x"0107",x"0289",
    x"03B9",x"00FF",x"0224",x"0046",x"01ED",x"0079",x"0209",x"0022",
    x"0275",x"0274",x"0271",x"0270",x"02A2",x"0042",x"0076",x"01DB",
    x"0057",x"02A1",x"0041",x"0071",x"0053",x"016B",x"020C",x"000B",
    x"0049",x"004E",x"0042",x"01CA",x"0242",x"031C",x"0004",x"0110",
    x"029B",x"0200",x"0003",x"0010",x"022C",x"0019",x"02B0",x"02B1",
    x"02B4",x"02B5",x"000D",x"0345",x"0104",x"022D",x"0071",x"0089",
    x"022C",x"002C",x"02B7",x"0275",x"0098",x"0004",x"0114",x"036C",
    x"0009",x"0288",x"0080",x"0224",x"007F",x"0281",x"031B",x"0009",
    x"028A",x"0342",x"0319",x"0204",x"01F3",x"02B7",x"0275",x"0004",
    x"0114",x"02F7",x"0229",x"008E",x"02B8",x"0001",x"0165",x"0206",
    x"002C",x"0048",x"0200",x"0029",x"0275",x"0004",x"0114",x"030F",
    x"0229",x"009C",x"02B8",x"0001",x"0165",x"0206",x"0006",x"0048",
    x"0200",x"0003",x"0275",x"02B8",x"0003",x"0270",x"008C",x"0098",
    x"0004",x"0114",x"036C",x"02F9",x"0003",x"0288",x"02BA",x"00FF",
    x"0040",x"0190",x"0011",x"0042",x"038A",x"01C2",x"00A1",x"02B0",
    x"0200",x"0003",x"0275",x"02B8",x"0003",x"0273",x"008C",x"02FC",
    x"0002",x"02F9",x"0004",x"028B",x"0004",x"0110",x"02FB",x"0043",
    x"0042",x"0004",x"0110",x"02FB",x"0043",x"0042",x"024B",x"0339",
    x"0004",x"02B3",x"02B7",x"0362",x"009B",x"0201",x"0008",x"0203",
    x"0008",x"0078",x"0209",x"0058",x"03BB",x"00FF",x"00AF",x"0223",
    x"0007",x"0060",x"00AF",x"0275",x"008D",x"0015",x"02AB",x"000D",
    x"02A9",x"0241",x"0319",x"0282",x"011C",x"0382",x"011A",x"02AA",
    x"0242",x"031A",x"02A8",x"0204",x"000C",x"0081",x"0082",x"03BA",
    x"00FF",x"01D1",x"0042",x"033D",x"000B",x"02E9",x"02EA",x"0200",
    x"0006",x"0053",x"0201",x"0003",x"0004",x"0114",x"0077",x"02A3",
    x"03BB",x"0300",x"0043",x"009D",x"0014",x"0001",x"02A3",x"0243",
    x"031C",x"0283",x"031B",x"02FB",x"0002",x"009C",x"0359",x"0261",
    x"020C",x"0004",x"0362",x"0224",x"011F",x"0014",x"0262",x"0015",
    x"022B",x"0124",x"020C",x"0011",x"0088",x"03C0",x"0319",x"0203",
    x"0007",x"0088",x"0050",x"0207",x"0003",x"0004",x"0110",x"03B1",
    x"0092",x"02B5",x"020B",x"005E",x"00AF",x"02BC",x"00FF",x"0041",
    x"01A1",x"0042",x"01A2",x"0015",x"0204",x"0031",x"0283",x"0319",
    x"0043",x"01A3",x"0343",x"0116",x"022E",x"0148",x"0343",x"0117",
    x"0225",x"014C",x"0283",x"031A",x"0043",x"01A3",x"0343",x"0118",
    x"022E",x"0154",x"0343",x"0119",x"0225",x"0158",x"01C0",x"0341",
    x"0116",x"020E",x"0005",x"0008",x"0341",x"0117",x"020D",x"0003",
    x"0004",x"0110",x"03C3",x"02B8",x"0002",x"0342",x"0118",x"020E",
    x"0033",x"0008",x"0342",x"0119",x"0205",x"002E",x"02B7",x"0379",
    x"00A7",x"0206",x"0009",x"01C0",x"0379",x"00B3",x"0205",x"0001",
    x"0008",x"0004",x"0110",x"03C3",x"037A",x"0067",x"0226",x"0182",
    x"02B8",x"0002",x"037A",x"0073",x"0205",x"0016",x"0008",x"0200",
    x"0013",x"0051",x"0030",x"0071",x"0038",x"01C0",x"0209",x"000B",
    x"0200",x"0008",x"0056",x"0030",x"0076",x"0038",x"02B8",x"0002",
    x"020A",x"0001",x"0008",x"0275",x"02BD",x"0001",x"0168",x"0206",
    x"0001",x"00ED",x"0271",x"0272",x"0281",x"031B",x"0009",x"00E9",
    x"02FD",x"0318",x"02AA",x"028B",x"024A",x"0082",x"0004",x"0114",
    x"00A1",x"02B2",x"02B1",x"02B7",x"0280",x"011C",x"0284",x"031B",
    x"0275",x"02FC",x"0002",x"02A3",x"02A5",x"0281",x"011A",x"0181",
    x"0224",x"01C4",x"0060",x"02A1",x"008A",x"03BA",x"00FF",x"01D1",
    x"0042",x"010B",x"0115",x"033C",x"000B",x"0263",x"0265",x"0220",
    x"0013",x"02F9",x"0005",x"028B",x"033B",x"0001",x"0225",x"00A3",
    x"024B",x"0280",x"011B",x"0204",x"0091",x"03BB",x"000F",x"022C",
    x"00AC",x"02BA",x"013B",x"00C2",x"03D3",x"0224",x"00B2",x"0009",
    x"028A",x"0004",x"0318",x"01B9",x"0280",x"0111",x"0064",x"02F8",
    x"0002",x"01C9",x"0200",x"0007",x"02B9",x"0001",x"0378",x"0003",
    x"020E",x"0001",x"0049",x"0275",x"0271",x"03B8",x"0006",x"0004",
    x"0114",x"003F",x"0273",x"0271",x"0008",x"0004",x"0114",x"003F",
    x"0010",x"0079",x"0050",x"02B1",x"0079",x"0050",x"02B2",x"02B1",
    x"02BD",x"0111",x"0268",x"026A",x"026B",x"0269",x"02B7",x"0275",
    x"01DB",x"0340",x"0104",x"022D",x"021F",x"0004",x"0114",x"036C",
    x"028C",x"0009",x"028A",x"0092",x"0224",x"0228",x"02F9",x"0004",
    x"02FA",x"0004",x"028B",x"006F",x"03BB",x"00FC",x"037B",x"00FC",
    x"0204",x"0005",x"0043",x"02CB",x"0209",x"000A",x"000F",x"028B",
    x"000B",x"009D",x"03BD",x"000F",x"0355",x"020C",x"0001",x"01EB",
    x"024B",x"03BB",x"000F",x"0006",x"03BC",x"0040",x"0204",x"0002",
    x"004B",x"0007",x"0051",x"000A",x"02D3",x"000B",x"02B7",x"0272",
    x"0082",x"0204",x"0019",x"03BA",x"00FF",x"01D0",x"0042",x"02C7",
    x"0115",x"006C",x"006E",x"006C",x"006E",x"006C",x"00C1",x"006E",
    x"02F2",x"00AF",x"006C",x"006E",x"0034",x"006C",x"006E",x"006C",
    x"006E",x"0068",x"00C1",x"006A",x"02F2",x"00AF",x"0275",x"02FC",
    x"0002",x"0001",x"02A1",x"0241",x"031C",x"0004",x"0118",x"018D",
    x"02B5",x"0281",x"031B",x"0009",x"028C",x"0011",x"00A4",x"0224",
    x"014C",x"0284",x"031C",x"00A4",x"0224",x"0151",x"0280",x"011B",
    x"00A7",x"0274",x"02BC",x"0019",x"0244",x"011E",x"02B7",x"02B9",
    x"00FF",x"0290",x"0040",x"03D8",x"0018",x"022C",x"0007",x"0011",
    x"022C",x"0008",x"00AF",x"0275",x"0270",x"0271",x"02BA",x"01FE",
    x"02BB",x"01FF",x"0004",x"0114",x"00B7",x"0008",x"0004",x"0114",
    x"027D",x"0290",x"0040",x"03D8",x"0018",x"0224",x"0009",x"02B8",
    x"01FF",x"0010",x"022C",x"0002",x"0290",x"0040",x"03D8",x"0018",
    x"0270",x"0004",x"0114",x"00B7",x"02B5",x"02B1",x"02B0",x"0220",
    x"0036",x"0001",x"03FF",x"03FE",x"0006",x"03FD",x"0004",x"0008",
    x"0000",x"0275",x"02B9",x"005A",x"0341",x"01FE",x"0204",x"000F",
    x"0341",x"01FF",x"0204",x"000B",x"02BC",x"011D",x"00A5",x"0001",
    x"02A0",x"0010",x"0268",x"0040",x"0268",x"020C",x"001C",x"02B8",
    x"0080",x"0240",x"0102",x"02BC",x"01FB",x"00A5",x"01DB",x"02A0",
    x"026B",x"02A1",x"026B",x"02A2",x"026B",x"0272",x"0004",x"0114",
    x"00C3",x"02B2",x"02BD",x"01FB",x"0268",x"0269",x"026A",x"02B8",
    x"00A0",x"0240",x"0102",x"02B9",x"011F",x"0282",x"01FF",x"0004",
    x"0114",x"012F",x"02B9",x"0120",x"0282",x"01FE",x"000F",x"0275",
    x"03FA",x"00FF",x"01C0",x"008B",x"02FB",x"0004",x"035A",x"025A",
    x"020C",x"0011",x"0093",x"03BB",x"001F",x"0066",x"0066",x"0062",
    x"00FA",x"033A",x"0058",x"0290",x"0004",x"0114",x"0268",x"0378",
    x"0001",x"020E",x"001D",x"008A",x"02FA",x"0002",x"0294",x"00A4",
    x"0204",x"000F",x"0270",x"0271",x"0273",x"01C0",x"0250",x"0010",
    x"00E4",x"02FC",x"0002",x"0004",x"0114",x"01EB",x"02B3",x"02B1",
    x"02B0",x"0084",x"0204",x"0048",x"020B",x"0055",x"0200",x"0028",
    x"0273",x"0271",x"0084",x"0338",x"0002",x"0060",x"02F9",x"0002",
    x"02C4",x"035D",x"0348",x"0248",x"0001",x"02A2",x"0204",x"0010",
    x"0004",x"0110",x"00AB",x"000C",x"00AB",x"0067",x"007B",x"0010",
    x"022C",x"0003",x"0004",x"0114",x"0205",x"02B8",x"0001",x"000F",
    x"01C0",x"02B1",x"0271",x"0004",x"0114",x"01EF",x"02B1",x"02B3",
    x"02B8",x"000F",x"01E4",x"0004",x"0114",x"01A6",x"0012",x"0013",
    x"0003",x"0001",x"0011",x"0019",x"0009",x"0008",x"0018",x"001C",
    x"000C",x"0004",x"0014",x"0016",x"0006",x"0002",x"036B",x"0204",
    x"0033",x"0010",x"0223",x"0005",x"0288",x"0082",x"03BA",x"00BF",
    x"03FA",x"0040",x"024A",x"03B8",x"00C0",x"022C",x"0100",x"0010",
    x"01E4",x"0200",x"002F",x"000C",x"009D",x"03BB",x"000F",x"0224",
    x"0014",x"01DD",x"022C",x"0017",x"02FC",x"0003",x"007B",x"0229",
    x"0004",x"022C",x"001E",x"00A0",x"0378",x"000B",x"0204",x"0004",
    x"020B",x"0004",x"02F8",x"000A",x"0338",x"000B",x"03B8",x"007F",
    x"03F8",x"0080",x"02BC",x"0002",x"0348",x"0224",x"0128",x"0248",
    x"0271",x"0274",x"0004",x"0114",x"01F9",x"02B4",x"02B1",x"0288",
    x"03B8",x"007F",x"02B5",x"02C4",x"035D",x"0001",x"02A2",x"0004",
    x"0014",x"00B1",x"0092",x"020C",x"0001",x"00AF",x"0339",x"011F",
    x"0097",x"0275",x"0004",x"0110",x"00AB",x"000C",x"00A9",x"02B5",
    x"0079",x"0044",x"0203",x"0001",x"0079",x"0229",x"0011",x"0004",
    x"001C",x"02AD",x"0275",x"0004",x"0118",x"03BB",x"03E9",x"0005",
    x"000C",x"0080",x"002B",x"0040",x"0018",x"000B",x"012B",x"03CF",
    x"0000",x"0018",x"002D",x"003B",x"0040",x"003B",x"002D",x"0018",
    x"0000",x"03E8",x"03D3",x"03C5",x"03C0",x"03C5",x"03D3",x"03E8",
    x"02A8",x"0275",x"0272",x"0004",x"0114",x"0237",x"0272",x"0004",
    x"0114",x"023D",x"02B0",x"0091",x"02B2",x"0200",x"0119",x"0275",
    x"0271",x"02F9",x"0004",x"0200",x"0004",x"0275",x"0271",x"02F9",
    x"0008",x"0270",x"0080",x"0203",x"0003",x"02F9",x"0008",x"0020",
    x"03B9",x"000F",x"0001",x"02F9",x"0018",x"0016",x"0289",x"0041",
    x"006D",x"006D",x"01D2",x"006D",x"006D",x"0078",x"0209",x"0001",
    x"00CA",x"0049",x"0080",x"022C",x"0007",x"004E",x"004A",x"02FA",
    x"0080",x"006E",x"006E",x"006E",x"006E",x"02B0",x"02B1",x"02B7",
    x"0040",x"0275",x"006C",x"0034",x"006C",x"006C",x"006C",x"02B7",
    x"0368",x"0205",x"0006",x"0368",x"0206",x"0002",x"0015",x"02A8",
    x"00AF",x"0015",x"02A8",x"000D",x"00AF",x"0275",x"0085",x"0204",
    x"0153",x"0271",x"0272",x"01D2",x"0280",x"035E",x"004C",x"004C",
    x"0081",x"03C0",x"035E",x"0041",x"0049",x"01C8",x"004D",x"01C8",
    x"0050",x"0280",x"035E",x"0050",x"0240",x"035E",x"0007",x"0052",
    x"0015",x"022C",x"0014",x"0190",x"0200",x"0134",x"0275",x"0271",
    x"0272",x"0081",x"0204",x"012E",x"01D2",x"000A",x"0060",x"022C",
    x"0003",x"0090",x"0004",x"0114",x"027D",x"0148",x"022D",x"0006",
    x"0200",x"0120",x"02B8",x"0001",x"0275",x"0004",x"0114",x"03C1",
    x"008C",x"0095",x"0082",x"00A9",x"0004",x"0118",x"0192",x"0004",
    x"0114",x"02D5",x"008D",x"02BB",x"0008",x"0001",x"02A1",x"0269",
    x"0013",x"022C",x"0005",x"0012",x"022C",x"0012",x"02B7",x"0275",
    x"0004",x"0114",x"02E6",x"011A",x"02B7",x"0275",x"0004",x"0114",
    x"02DB",x"011A",x"02B7",x"0270",x"0271",x"02A9",x"0275",x"0004",
    x"0114",x"0345",x"0018",x"0388",x"0200",x"000B",x"0270",x"0271",
    x"02A9",x"0275",x"0004",x"0114",x"0345",x"0085",x"0018",x"0388",
    x"01E8",x"0248",x"02B5",x"02B1",x"02B0",x"0275",x"02B7",x"0275",
    x"0272",x"0004",x"0114",x"0377",x"02B5",x"0275",x"00A8",x"03BD",
    x"00FF",x"01E8",x"0040",x"0102",x"0203",x"0001",x"0022",x"012B",
    x"0203",x"0001",x"0023",x"02B0",x"0271",x"0200",x"0013",x"0275",
    x"0098",x"0004",x"0114",x"0377",x"0271",x"0272",x"0273",x"0004",
    x"0114",x"0372",x"0333",x"0203",x"0001",x"0023",x"0332",x"0203",
    x"0001",x"0022",x"00A1",x"03BC",x"00FF",x"01E1",x"0041",x"0111",
    x"0209",x"0001",x"011C",x"008D",x"02B1",x"0082",x"0083",x"02B7",
    x"0275",x"008D",x"02A1",x"0269",x"0010",x"022C",x"0004",x"02B7",
    x"0275",x"01ED",x"0270",x"0265",x"0010",x"022C",x"0003",x"02B0",
    x"02B7",x"0275",x"008D",x"0220",x"000A",x"0275",x"0085",x"02B8",
    x"0001",x"000F",x"0048",x"0015",x"0223",x"0003",x"02B7",x"0275",
    x"03B8",x"00FF",x"0040",x"03B9",x"00FF",x"01C8",x"02B7",x"0275",
    x"0270",x"0004",x"0114",x"0268",x"0081",x"02B0",x"0220",x"00F5",
    x"0275",x"0009",x"0288",x"0011",x"0080",x"02B7",x"0088",x"0338",
    x"031D",x"0064",x"0060",x"00AF",x"0081",x"004D",x"0049",x"02F9",
    x"031D",x"00AF",x"0275",x"0004",x"0114",x"036C",x"000F",x"0275",
    x"008D",x"02FD",x"0002",x"02AA",x"0042",x"03BA",x"00FF",x"02AB",
    x"0043",x"03BB",x"00FF",x"02B7",x"02A0",x"0040",x"03B8",x"00FF",
    x"02A1",x"0041",x"03B9",x"00FF",x"0275",x"0270",x"0110",x"0020",
    x"0270",x"0271",x"0004",x"011C",x"01DB",x"02B0",x"0084",x"0118",
    x"0020",x"0270",x"0272",x"0004",x"011C",x"01DB",x"02F2",x"02B1",
    x"02B0",x"02B3",x"02B7",x"0275",x"0004",x"0114",x"0384",x"0083",
    x"008C",x"0091",x"02B5",x"0004",x"031C",x"0223",x"0009",x"01C0",
    x"0248",x"0011",x"00AF",x"0275",x"02BA",x"0007",x"0090",x"0004",
    x"0114",x"036C",x"0004",x"0114",x"03AE",x"0012",x"0223",x"0009",
    x"02B7",x"0271",x"0272",x"0273",x"0274",x"0001",x"02BC",x"00D0",
    x"0017",x"0274",x"0275",x"00B5",x"033D",x"0003",x"02AC",x"02B7",
    x"02B4",x"02B3",x"02B2",x"02B1",x"02B7",x"0275",x"0004",x"0110",
    x"00AB",x"0002",x"02BC",x"0125",x"0001",x"02A8",x"0001",x"02AB",
    x"0080",x"0204",x"003A",x"00A2",x"0001",x"02A1",x"0339",x"0001",
    x"0225",x"000D",x"0094",x"0261",x"0041",x"0261",x"022C",x"0013",
    x"0094",x"0263",x"0043",x"0263",x"0275",x"00BD",x"02FD",x"0004",
    x"0274",x"0087",x"02B4",x"02B5",x"0220",x"0021",x"0275",x"0004",
    x"0110",x"00AB",x"0002",x"02BC",x"0125",x"0001",x"02A8",x"0080",
    x"0204",x"0013",x"0001",x"02A8",x"0260",x"0040",x"0260",x"0220",
    x"000B",x"0275",x"0274",x"0004",x"0110",x"00AB",x"0002",x"02B4",
    x"0129",x"0069",x"02F9",x"0125",x"008D",x"02B7",x"0275",x"0271",
    x"0272",x"008D",x"0001",x"02A8",x"0001",x"02AA",x"004A",x"0062",
    x"0004",x"0118",x"0011",x"026A",x"0042",x"026A",x"02B2",x"02B1",
    x"02B7",x"0275",x"0271",x"0004",x"0118",x"0011",x"0200",x"0015",
    x"0275",x"0271",x"0004",x"0118",x"0011",x"0001",x"02A8",x"0048",
    x"0007",x"0070",x"0200",x"0009",x"0275",x"0271",x"0004",x"0118",
    x"0011",x"0001",x"02A8",x"0048",x"0060",x"0248",x"0009",x"0040",
    x"0248",x"02B1",x"02B7",x"0275",x"0271",x"0274",x"009D",x"0265",
    x"0281",x"0105",x"0071",x"0201",x"0004",x"0001",x"03BD",x"00FF",
    x"00DF",x"0010",x"022C",x"000C",x"02B4",x"02B1",x"02B7",x"0275",
    x"0007",x"008D",x"0200",x"0010",x"0275",x"0007",x"008D",x"0200",
    x"0001",x"0006",x"004B",x"0073",x"0275",x"0004",x"0118",x"0053",
    x"02B5",x"0200",x"0003",x"0006",x"004B",x"0073",x"0273",x"02A8",
    x"03B8",x"007F",x"020C",x"0005",x"009B",x"02B3",x"020B",x"0076",
    x"00AF",x"0338",x"0020",x"004C",x"0048",x"01D8",x"0260",x"0280",
    x"0105",x"0070",x"0221",x"0014",x"0001",x"03BB",x"00FF",x"00DF",
    x"0220",x"001A",x"0001",x"000A",x"0064",x"03E8",x"0275",x"0270",
    x"0088",x"0004",x"0118",x"0053",x"02B0",x"0004",x"0114",x"03C1",
    x"004B",x"0007",x"0073",x"0200",x"001C",x"0275",x"0004",x"0114",
    x"03C1",x"02BA",x"0080",x"01DA",x"0200",x"0014",x"0275",x"0270",
    x"0280",x"0105",x"0070",x"0201",x"0006",x"0001",x"02BD",x"00FF",
    x"00DF",x"01AB",x"01AA",x"02B0",x"02B7",x"0275",x"0004",x"0114",
    x"03C1",x"009A",x"0080",x"0203",x"0009",x"0020",x"0011",x"02BD",
    x"0068",x"01DD",x"0265",x"0004",x"0118",x"00B6",x"00F9",x"0339",
    x"003E",x"028D",x"0168",x"0203",x"000D",x"0015",x"0204",x"000A",
    x"009B",x"020B",x"0004",x"0262",x"0004",x"0118",x"00B6",x"0011",
    x"0220",x"0010",x"02BA",x"0080",x"0308",x"020B",x"0004",x"02FA",
    x"0008",x"0220",x"0006",x"02C8",x"01DA",x"0262",x"0004",x"0118",
    x"00B6",x"028A",x"0011",x"0012",x"022C",x"0013",x"02B7",x"0004",
    x"0018",x"0110",x"0000",x"0000",x"004C",x"0019",x"0000",x"0000",
    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
    x"0244",x"035D",x"02BC",x"0131",x"0262",x"0339",x"0200",x"0261",
    x"0260",x"02FC",x"0003",x"0265",x"00A8",x"0040",x"0260",x"0263",
    x"0043",x"0263",x"02BC",x"0132",x"02A1",x"02F9",x"0200",x"02A0",
    x"01ED",x"0265",x"0265",x"0265",x"02FC",x"0002",x"0001",x"03E5",
    x"024D",x"0011",x"0010",x"022C",x"0004",x"02B7",x"0275",x"0280",
    x"0149",x"0080",x"0224",x"003D",x"0280",x"035F",x"0001",x"0338",
    x"000A",x"0016",x"022B",x"0045",x"0378",x"0014",x"022E",x"0049",
    x"0004",x"011C",x"02BD",x"02B7",x"0275",x"0341",x"0131",x"022C",
    x"0052",x"0378",x"000A",x"0224",x"0032",x"02BD",x"0134",x"02AA",
    x"0378",x"000B",x"020C",x"000B",x"00B8",x"0338",x"0057",x"0283",
    x"035D",x"0240",x"035D",x"0001",x"02A8",x"0001",x"02AF",x"02BD",
    x"0133",x"036A",x"0224",x"0034",x"000A",x"026A",x"00AC",x"0001",
    x"02A9",x"0049",x"0271",x"004D",x"02F1",x"00C1",x"0261",x"0041",
    x"0261",x"0281",x"0132",x"02F9",x"0200",x"004C",x"0048",x"02F8",
    x"0080",x"02FD",x"0002",x"0001",x"03E8",x"028B",x"0248",x"0098",
    x"0011",x"0012",x"022C",x"0006",x"02B7",x"0275",x"0004",x"0114",
    x"036C",x"000F",x"0275",x"0004",x"0114",x"0366",x"0271",x"02F9",
    x"0006",x"01ED",x"024D",x"0081",x"02F9",x"013B",x"024D",x"02B1",
    x"02B7",x"0007",x"000F",x"0006",x"0053",x"0275",x"0200",x"0019",
    x"0275",x"0004",x"0114",x"0366",x"000F",x"0275",x"0004",x"0114",
    x"036C",x"0085",x"02FD",x"013B",x"026B",x"02F9",x"0007",x"024A",
    x"02B5",x"0007",x"000F",x"0006",x"0275",x"0053",x"0004",x"0114",
    x"036C",x"0004",x"0114",x"03C1",x"02F9",x"0002",x"008C",x"0274",
    x"0273",x"0093",x"03BB",x"00FF",x"01DA",x"0042",x"0004",x"0114",
    x"03A3",x"02B1",x"0098",x"0203",x"0001",x"0023",x"00DB",x"0079",
    x"0049",x"0053",x"0273",x"0271",x"0093",x"0004",x"011C",x"01DC",
    x"02B1",x"02B5",x"00A0",x"0203",x"0001",x"0024",x"00E4",x"00E4",
    x"016C",x"0205",x"0005",x"03BD",x"0001",x"01E5",x"03FD",x"0002",
    x"0275",x"0094",x"0004",x"011C",x"01DC",x"0091",x"009A",x"0004",
    x"011C",x"01F8",x"009A",x"0083",x"00A1",x"0004",x"011C",x"01F8",
    x"03BB",x"00FF",x"03B8",x"00FF",x"0040",x"01D8",x"02B3",x"02B4",
    x"02FC",x"0002",x"0260",x"007B",x"0229",x"006D",x"01C9",x"01D2",
    x"0004",x"0114",x"0077",x"007B",x"0201",x"0001",x"008A",x"0092",
    x"0203",x"0001",x"0022",x"0099",x"0041",x"0061",x"0062",x"0004",
    x"011C",x"01F8",x"0080",x"020C",x"0003",x"0014",x"0260",x"0008",
    x"000C",x"0260",x"00A1",x"0004",x"0114",x"0366",x"02B7",x"0275",
    x"0272",x"01ED",x"0021",x"020D",x"0004",x"02FD",x"0008",x"0020",
    x"0021",x"0080",x"020D",x"0006",x"008A",x"0020",x"0081",x"0090",
    x"02FD",x"0004",x"008A",x"004E",x"0150",x"020E",x"0012",x"000D",
    x"0082",x"010A",x"004E",x"0150",x"0206",x"000B",x"000D",x"0022",
    x"0151",x"020E",x"0006",x"000D",x"004C",x"0141",x"0206",x"0001",
    x"000D",x"00A9",x"03B9",x"000F",x"02B2",x"02B7",x"0275",x"008D",
    x"000F",x"02A8",x"0245",x"0143",x"00A9",x"0041",x"0241",x"0144",
    x"0004",x"0110",x"00AB",x"0002",x"00A9",x"02B5",x"0004",x"0318",
    x"0031",x"0275",x"02BD",x"0143",x"0001",x"02AF",x"0343",x"0146",
    x"0205",x"0019",x"020E",x"0004",x"0073",x"0201",x"0014",x"0053",
    x"0243",x"0146",x"00A7",x"0275",x"0270",x"0271",x"02BC",x"01F0",
    x"02B8",x"000E",x"0004",x"0114",x"0338",x"02B8",x"0038",x"0240",
    x"01F8",x"02B1",x"02B0",x"02B7",x"02BC",x"0002",x"0244",x"0148",
    x"0245",x"035F",x"0004",x"0118",x"0283",x"0240",x"0149",x"01C0",
    x"0240",x"0145",x"02B7",x"033E",x"0003",x"0004",x"0118",x"0283",
    x"02B8",x"00FF",x"0240",x"0145",x"02B7",x"0280",x"0145",x"0010",
    x"020B",x"000A",x"0275",x"01C0",x"0240",x"0145",x"0240",x"0149",
    x"0240",x"0146",x"0287",x"035F",x"00AF",x"02B9",x"0148",x"0288",
    x"0010",x"0248",x"022C",x"0007",x"0282",x"0147",x"024A",x"03C0",
    x"0145",x"022C",x"000E",x"0275",x"02C7",x"0149",x"0248",x"02B7",
    x"0200",x"0059",x"0200",x"007E",x"0200",x"008B",x"0200",x"009A",
    x"0200",x"00BF",x"0200",x"0122",x"005D",x"000D",x"009C",x"000C",
    x"00E7",x"000B",x"003C",x"000B",x"009B",x"000A",x"0003",x"000A",
    x"0072",x"0009",x"00EB",x"0008",x"006B",x"0008",x"00F2",x"0007",
    x"007F",x"0007",x"0014",x"0007",x"0275",x"0273",x"0274",x"01C9",
    x"0285",x"035F",x"02AB",x"0245",x"035F",x"009B",x"0224",x"005C",
    x"007F",x"0055",x"007B",x"0051",x"01D2",x"007B",x"0052",x"037B",
    x"003F",x"0224",x"0012",x"0009",x"004D",x"0098",x"0204",x"0014",
    x"01E4",x"02BD",x"000C",x"000C",x"012B",x"0223",x"0003",x"00DD",
    x"00ED",x"00FD",x"033D",x"003E",x"0001",x"02A8",x"0060",x"0014",
    x"022C",x"0003",x"0008",x"0060",x"02B4",x"02B3",x"02B7",x"02B8",
    x"0002",x"0220",x"0096",x"0004",x"0118",x"02F4",x"0092",x"0204",
    x"0006",x"0339",x"0002",x"02BD",x"0004",x"0245",x"0149",x"0004",
    x"0118",x"03AE",x"02BD",x"01F0",x"0268",x"0268",x"0268",x"01D2",
    x"026A",x"0040",x"0268",x"0268",x"0268",x"01D2",x"026A",x"02FD",
    x"0003",x"0080",x"0204",x"0002",x"02B8",x"000F",x"0268",x"0268",
    x"0268",x"02B7",x"0004",x"0118",x"0283",x"02B9",x"0002",x"0004",
    x"0118",x"03AE",x"0241",x"0149",x"02B7",x"02B8",x"0006",x"0220",
    x"00CC",x"0004",x"0118",x"02F4",x"0092",x"0204",x"0006",x"0339",
    x"0002",x"02BD",x"0008",x"0245",x"0149",x"0004",x"0118",x"037F",
    x"0220",x"002C",x"0004",x"0118",x"0283",x"02B9",x"0002",x"0004",
    x"0118",x"03AE",x"02B9",x"0006",x"0241",x"0149",x"02B7",x"0275",
    x"0004",x"0118",x"03AE",x"02BD",x"01F0",x"0268",x"0060",x"0268",
    x"0060",x"0268",x"01D2",x"026A",x"004C",x"0040",x"0268",x"0034",
    x"0060",x"0268",x"0060",x"0268",x"02B7",x"02B8",x"000A",x"0220",
    x"0104",x"0004",x"0118",x"02F4",x"0004",x"0118",x"037F",x"02B9",
    x"0020",x"0269",x"02FD",x"0002",x"026A",x"0080",x"0204",x"0002",
    x"02B8",x"003F",x"0268",x"0268",x"0268",x"02B7",x"0275",x"0270",
    x"0285",x"0147",x"01C0",x"00C8",x"0015",x"022C",x"0003",x"0240",
    x"0148",x"02B0",x"02B7",x"02BB",x"0080",x"000F",x"02AB",x"0004",
    x"0018",x"0276",x"02BC",x"0002",x"0244",x"0148",x"0245",x"035F",
    x"0014",x"0240",x"0159",x"0244",x"014A",x"02B8",x"000A",x"02BC",
    x"014B",x"0004",x"0114",x"0338",x"02B8",x"000C",x"0220",x"013A",
    x"0000",x"0002",x"0004",x"000B",x"001A",x"003B",x"0078",x"00F5",
    x"0007",x"0000",x"0007",x"0009",x"000C",x"0012",x"0013",x"0000",
    x"0110",x"002F",x"00A4",x"00E8",x"00C4",x"0137",x"014D",x"016E",
    x"00C1",x"0143",x"0043",x"0076",x"00CF",x"00DD",x"0162",x"00B0",
    x"0127",x"00CB",x"0142",x"013C",x"0129",x"0123",x"02BB",x"01F0",
    x"02BC",x"014B",x"02A0",x"02A1",x"00C8",x"0021",x"0014",x"0261",
    x"0004",x"0114",x"0268",x"0204",x"0008",x"02D8",x"0258",x"009A",
    x"02FA",x"0004",x"0040",x"02D0",x"0250",x"000B",x"037C",x"0151",
    x"022C",x"0017",x"02BA",x"0155",x"02A0",x"0004",x"0114",x"0268",
    x"02D0",x"0004",x"0114",x"0270",x"0004",x"007F",x"0250",x"0064",
    x"02FB",x"0006",x"0258",x"000B",x"000A",x"000B",x"02A0",x"0080",
    x"0204",x"0007",x"02D0",x"0250",x"0064",x"0060",x"03B8",x"000F",
    x"0258",x"037C",x"0155",x"022C",x"0010",x"0280",x"014A",x"0010",
    x"0240",x"014A",x"022C",x"01B0",x"0284",x"035F",x"00BD",x"0015",
    x"0275",x"02A0",x"01C9",x"033D",x"006E",x"00AA",x"02FA",x"0006",
    x"000A",x"0078",x"0051",x"0369",x"022D",x"0005",x"033D",x"0002",
    x"0329",x"0015",x"0329",x"02D2",x"00CA",x"02BB",x"01F0",x"02D7",
    x"01D2",x"007C",x"0056",x"02A1",x"00D3",x"0259",x"02FB",x"0004",
    x"004D",x"004D",x"004D",x"005D",x"0054",x"0081",x"0065",x"0065",
    x"0258",x"037A",x"0003",x"0204",x"0014",x"01C0",x"0095",x"00ED",
    x"02FD",x"014B",x"0268",x"0268",x"0088",x"0224",x"01EB",x"0113",
    x"02FB",x"0007",x"0011",x"020C",x"00C8",x"02B8",x"0030",x"0200",
    x"00C4",x"02FB",x"0003",x"0298",x"0258",x"0258",x"02B7",x"02A1",
    x"01D2",x"007D",x"0056",x"02BD",x"014B",x"037A",x"0003",x"020C",
    x"0005",x"0269",x"0268",x"0269",x"0268",x"01D2",x"00D5",x"00D5",
    x"0269",x"0268",x"02B7",x"0004",x"011C",x"00C2",x"029D",x"02FB",
    x"0004",x"0299",x"03B9",x"000F",x"0041",x"01E9",x"0004",x"011C",
    x"00EC",x"0041",x"0259",x"033B",x"0004",x"0041",x"0259",x"000B",
    x"037B",x"01F3",x"022C",x"0015",x"02B7",x"0041",x"006D",x"006D",
    x"006D",x"006D",x"0008",x"00C0",x"0245",x"035F",x"0082",x"0090",
    x"01ED",x"000D",x"0060",x"022C",x"0003",x"00A8",x"0004",x"0114",
    x"027D",x"0150",x"022D",x"000C",x"0287",x"035F",x"0004",x"011C",
    x"00C2",x"02BB",x"014B",x"0299",x"0041",x"006D",x"006D",x"006D",
    x"006D",x"0004",x"011C",x"00EC",x"0259",x"02FB",x"0002",x"037B",
    x"0151",x"022C",x"000F",x"02B7",x"0275",x"0082",x"008D",x"01C9",
    x"007A",x"0209",x"0003",x"0025",x"000F",x"00E9",x"0012",x"0223",
    x"0003",x"0082",x"007A",x"0209",x"0001",x"0025",x"006D",x"006D",
    x"0009",x"0069",x"00E9",x"02B7",x"02FB",x"0008",x"0258",x"0081",
    x"0065",x"0061",x"0188",x"01C9",x"02FB",x"0002",x"0200",x"0004",
    x"02FB",x"000A",x"02B9",x"0030",x"02BA",x"0151",x"01ED",x"000A",
    x"000B",x"0078",x"0209",x"0002",x"0259",x"0255",x"022C",x"0008",
    x"02B7",x"0240",x"01FA",x"02B7",x"0240",x"01F9",x"004C",x"0240",
    x"0155",x"01C0",x"000F",x"02A0",x"0240",x"0151",x"02B7",x"0281",
    x"0155",x"0004",x"011C",x"00C2",x"0004",x"011C",x"00EC",x"0241",
    x"0155",x"0065",x"0241",x"01F9",x"02B7",x"0281",x"0151",x"0004",
    x"011C",x"00BD",x"0004",x"011C",x"00EC",x"0241",x"0151",x"02B7",
    x"02FB",x"000B",x"01D2",x"007C",x"0056",x"01C9",x"037A",x"0003",
    x"020C",x"0002",x"0009",x"01D2",x"00D3",x"009D",x"0268",x"0089",
    x"0204",x"0002",x"0268",x"0268",x"02BD",x"0156",x"00D5",x"004C",
    x"0048",x"02FA",x"0152",x"01DB",x"0268",x"0253",x"0089",x"0224",
    x"02D5",x"0268",x"0268",x"000A",x"0253",x"000A",x"0253",x"02B7",
    x"01D2",x"007C",x"0056",x"0040",x"02BD",x"0152",x"004C",x"006C",
    x"0040",x"037A",x"0003",x"020C",x"0003",x"0268",x"0268",x"000F",
    x"00D5",x"0268",x"02B7",x"0008",x"0240",x"0147",x"02B7",x"0001",
    x"02A7",x"02B5",x"0074",x"020A",x"0004",x"0001",x"02BC",x"0093",
    x"001A",x"0244",x"035F",x"0229",x"02EF",x"0220",x"02EE",x"01DB",
    x"007C",x"0057",x"0200",x"0002",x"0083",x"02A0",x"02FB",x"0159",
    x"0258",x"02B7",x"02A0",x"0008",x"0080",x"0224",x"0313",x"0240",
    x"014A",x"0244",x"035F",x"02B5",x"02B7",x"02A1",x"01D2",x"007D",
    x"0056",x"02FA",x"0159",x"0295",x"0015",x"020B",x"0003",x"0255",
    x"0224",x"0015",x"0041",x"006D",x"006D",x"006D",x"006D",x"00CC",
    x"0220",x"001D",x"02A1",x"007D",x"0054",x"0079",x"0050",x"0008",
    x"0004",x"011C",x"00C4",x"00C8",x"0220",x"0029",x"02A1",x"01DB",
    x"007D",x"0057",x"007D",x"0054",x"0008",x"0004",x"011C",x"00C4",
    x"00C8",x"0220",x"003C",x"0081",x"0273",x"01DB",x"01D2",x"0080",
    x"0203",x"0002",x"0020",x"000B",x"0089",x"0203",x"0002",x"0021",
    x"000B",x"0200",x"0002",x"00C2",x"0048",x"0079",x"0221",x"0004",
    x"022C",x"0005",x"007B",x"0209",x"0001",x"0022",x"02B3",x"00AF",
    x"0090",x"0078",x"00C1",x"0273",x"01C0",x"02BB",x"0001",x"0092",
    x"0204",x"001F",x"0203",x"0002",x"0022",x"0008",x"000F",x"004B",
    x"005A",x"0229",x"0003",x"0072",x"0089",x"0203",x"0002",x"0021",
    x"0008",x"0078",x"0073",x"01C0",x"0062",x"0151",x"0205",x"0002",
    x"0111",x"0007",x"0050",x"007B",x"0229",x"0009",x"0204",x"0001",
    x"0020",x"02B3",x"00AF",x"0275",x"008A",x"0062",x"0272",x"0271",
    x"0004",x"011C",x"01F8",x"02B1",x"02B2",x"00C2",x"0062",x"0110",
    x"0203",x"0001",x"0020",x"0378",x"0002",x"0223",x"0010",x"02B7",
    x"0275",x"02B8",x"00F0",x"02BC",x"0200",x"0004",x"0114",x"0338",
    x"02BC",x"0216",x"0001",x"02B8",x"002F",x"0005",x"0260",x"000C",
    x"037C",x"021E",x"020C",x"0003",x"000C",x"0338",x"0008",x"0010",
    x"037C",x"0227",x"022C",x"000D",x"02B8",x"0082",x"0240",x"0102",
    x"0002",x"0340",x"0102",x"0224",x"0003",x"02BB",x"0007",x"0004",
    x"0110",x"00AB",x"000A",x"0274",x"02A8",x"0275",x"02B9",x"0002",
    x"02BC",x"02D2",x"0004",x"0118",x"00C5",x"02B4",x"00A1",x"0001",
    x"02BA",x"002D",x"0005",x"0012",x"02A0",x"0080",x"022C",x"0004",
    x"0062",x"0094",x"0004",x"0118",x"0067",x"02B1",x"0289",x"0045",
    x"0203",x"0005",x"00AC",x"00BD",x"02FD",x"0003",x"00A7",x"0004",
    x"0115",x"00C3",x"0003",x"00A9",x"03B9",x"00FF",x"020C",x"0002",
    x"01E9",x"0041",x"008A",x"03B9",x"001F",x"0011",x"02B8",x"0003",
    x"020C",x"0010",x"0048",x"0066",x"0066",x"007E",x"0202",x"0008",
    x"0010",x"007A",x"0201",x"0004",x"0010",x"007A",x"0229",x"0012",
    x"022C",x"0014",x"0240",x"0103",x"02B7",x"0281",x"0149",x"0089",
    x"020C",x"0001",x"00A7",x"00AF",x"0275",x"0004",x"0118",x"03BE",
    x"00FF",x"02CF",x"0004",x"001C",x"02AD",x"02B8",x"0005",x"0200",
    x"0003",x"0004",x"001C",x"02AD",x"0275",x"0004",x"0118",x"03BB",
    x"0040",x"0018",x"0048",x"0030",x"0044",x"0060",x"000C",x"0033",
    x"0389",x"020B",x"00C3",x"03F8",x"02CF",x"0275",x"0004",x"0118",
    x"03BB",x"0279",x"03ED",x"0105",x"01A5",x"0062",x"006A",x"01EB",
    x"0002",x"000A",x"000F",x"03FF",x"008F",x"0013",x"000F",x"0000",
    x"0013",x"0019",x"0003",x"0061",x"02E9",x"0280",x"0050",x"015B",
    x"0001",x"03F8",x"03EB",x"0013",x"002E",x"0023",x"0016",x"0001",
    x"000C",x"016B",x"0001",x"03F4",x"00C3",x"03E6",x"0001",x"0008",
    x"03EB",x"02F9",x"0157",x"002E",x"0013",x"0019",x"0003",x"0025",
    x"02C9",x"0280",x"0200",x"0308",x"0240",x"03EB",x"02F9",x"0097",
    x"0040",x"0003",x"0354",x"03F2",x"03FA",x"000F",x"0002",x"008F",
    x"0027",x"03F9",x"03CF",x"02B8",x"000E",x"0275",x"0004",x"0118",
    x"03BB",x"0389",x"0340",x"0028",x"0348",x"0029",x"0344",x"002A",
    x"006B",x"02C0",x"0030",x"02F5",x"0023",x"03D0",x"02CF",x"0275",
    x"0004",x"0110",x"00AB",x"0008",x"000F",x"0274",x"0275",x"0001",
    x"02BB",x"00DF",x"0036",x"009C",x"02FC",x"003A",x"02BD",x"0200",
    x"0298",x"000B",x"02BA",x"0004",x"02A1",x"0041",x"007C",x"0075",
    x"0065",x"0065",x"0065",x"0269",x"0012",x"022C",x"000A",x"037D",
    x"02E7",x"0225",x"0012",x"02B5",x"02A8",x"00AB",x"0001",x"02BD",
    x"0000",x"0038",x"00B9",x"0011",x"0271",x"0299",x"000B",x"0079",
    x"01D2",x"0209",x"0002",x"029A",x"000B",x"0270",x"0275",x"0273",
    x"02BC",x"02E8",x"007A",x"0209",x"0002",x"02BF",x"0213",x"007A",
    x"0201",x"003F",x"007A",x"0209",x"0004",x"01DB",x"0042",x"02BF",
    x"0200",x"0004",x"0100",x"02D3",x"0001",x"02BC",x"0000",x"0030",
    x"007A",x"0201",x"000F",x"0004",x"0110",x"00AB",x"0006",x"00AC",
    x"0090",x"03B8",x"0002",x"0204",x"0005",x"01C2",x"0001",x"02BC",
    x"0000",x"0038",x"0041",x"004D",x"007E",x"0075",x"0041",x"0280",
    x"02E6",x"00C1",x"0102",x"0204",x"0006",x"02B2",x"033A",x"0002",
    x"0272",x"0082",x"000A",x"0242",x"02E6",x"004D",x"00C9",x"00CC",
    x"02B9",x"02E8",x"02B8",x"0008",x"0004",x"0114",x"0330",x"02BF",
    x"0247",x"0088",x"03B8",x"0080",x"01C1",x"007A",x"0050",x"01DB",
    x"007E",x"0057",x"007A",x"0053",x"0078",x"0052",x"004C",x"0040",
    x"009B",x"020C",x"0003",x"0083",x"004F",x"01C0",x"0270",x"0273",
    x"0004",x"0100",x"02C3",x"02B5",x"02B8",x"0200",x"0060",x"0015",
    x"0223",x"0003",x"0042",x"004D",x"01D1",x"03F1",x"004D",x"004D",
    x"0004",x"0100",x"02DC",x"0059",x"0229",x"0005",x"0059",x"0209",
    x"000D",x"0060",x"020C",x"0002",x"02B8",x"0100",x"0004",x"0100",
    x"02DC",x"0059",x"0229",x"000A",x"0220",x"0015",x"0048",x"03B8",
    x"01FF",x"020C",x"0001",x"0008",x"0004",x"0100",x"02DC",x"0059",
    x"0229",x"000B",x"0220",x"0023",x"0000",x"0000",x"0000",x"0000");

  CONSTANT INIT_GROM : arr8 := (
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"30",x"30",x"30",x"30",x"30",x"00",x"30",x"00",
    x"66",x"66",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"14",x"3E",x"14",x"3E",x"14",x"00",x"00",
    x"10",x"FE",x"D0",x"FE",x"16",x"D6",x"FE",x"10",x"00",x"62",x"64",x"08",x"10",x"26",x"46",x"00",
    x"10",x"7C",x"60",x"38",x"60",x"7C",x"10",x"00",x"10",x"20",x"40",x"00",x"00",x"00",x"00",x"00",
    x"0E",x"08",x"08",x"08",x"08",x"08",x"08",x"0E",x"70",x"10",x"10",x"10",x"10",x"10",x"10",x"70",
    x"10",x"38",x"6C",x"38",x"10",x"00",x"00",x"00",x"00",x"18",x"18",x"7E",x"18",x"18",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"08",x"00",x"00",x"00",x"7E",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"01",x"02",x"04",x"08",x"10",x"20",x"40",x"80",
    x"00",x"FE",x"C6",x"D6",x"D6",x"C6",x"FE",x"00",x"00",x"38",x"18",x"18",x"18",x"18",x"7E",x"00",
    x"00",x"7E",x"66",x"06",x"7E",x"60",x"7E",x"00",x"00",x"7E",x"06",x"3C",x"06",x"06",x"7E",x"00",
    x"00",x"66",x"66",x"66",x"7E",x"06",x"06",x"00",x"00",x"7E",x"60",x"7E",x"06",x"66",x"7E",x"00",
    x"00",x"7E",x"60",x"7E",x"66",x"66",x"7E",x"00",x"00",x"7E",x"06",x"0C",x"18",x"30",x"30",x"00",
    x"00",x"7E",x"66",x"3C",x"66",x"66",x"7E",x"00",x"00",x"7E",x"66",x"66",x"7E",x"06",x"7E",x"00",
    x"00",x"00",x"18",x"18",x"00",x"18",x"18",x"00",x"00",x"00",x"18",x"18",x"00",x"18",x"18",x"08",
    x"00",x"06",x"18",x"60",x"18",x"06",x"00",x"00",x"00",x"00",x"7E",x"00",x"7E",x"00",x"00",x"00",
    x"00",x"60",x"18",x"06",x"18",x"60",x"00",x"00",x"7E",x"66",x"06",x"1E",x"18",x"00",x"18",x"00",
    x"FE",x"82",x"BA",x"AA",x"BE",x"80",x"FE",x"00",x"7E",x"66",x"66",x"66",x"7E",x"66",x"66",x"00",
    x"7E",x"66",x"66",x"7C",x"66",x"66",x"7E",x"00",x"7E",x"66",x"60",x"60",x"60",x"66",x"7E",x"00",
    x"7C",x"66",x"66",x"66",x"66",x"66",x"7C",x"00",x"7E",x"60",x"60",x"7C",x"60",x"60",x"7E",x"00",
    x"7E",x"60",x"60",x"7C",x"60",x"60",x"60",x"00",x"7E",x"66",x"60",x"6E",x"66",x"66",x"7E",x"00",
    x"66",x"66",x"66",x"7E",x"66",x"66",x"66",x"00",x"7E",x"18",x"18",x"18",x"18",x"18",x"7E",x"00",
    x"06",x"06",x"06",x"06",x"66",x"66",x"7E",x"00",x"66",x"66",x"6C",x"78",x"66",x"66",x"66",x"00",
    x"60",x"60",x"60",x"60",x"60",x"60",x"7E",x"00",x"82",x"C6",x"EE",x"FE",x"D6",x"D6",x"C6",x"00",
    x"46",x"66",x"76",x"7E",x"6E",x"66",x"62",x"00",x"7E",x"66",x"66",x"66",x"66",x"66",x"7E",x"00",
    x"7E",x"66",x"66",x"66",x"7E",x"60",x"60",x"00",x"7E",x"66",x"66",x"66",x"66",x"6E",x"7E",x"03",
    x"7E",x"66",x"66",x"66",x"7C",x"66",x"66",x"00",x"7E",x"66",x"60",x"7E",x"06",x"66",x"7E",x"00",
    x"7E",x"18",x"18",x"18",x"18",x"18",x"18",x"00",x"66",x"66",x"66",x"66",x"66",x"66",x"7E",x"00",
    x"66",x"66",x"66",x"24",x"3C",x"18",x"18",x"00",x"C6",x"C6",x"D6",x"D6",x"FE",x"6C",x"6C",x"00",
    x"66",x"66",x"3C",x"18",x"3C",x"66",x"66",x"00",x"66",x"66",x"66",x"66",x"7E",x"18",x"18",x"00",
    x"7E",x"06",x"0C",x"18",x"30",x"60",x"7E",x"00",x"1E",x"18",x"18",x"18",x"18",x"18",x"18",x"1E",
    x"80",x"40",x"20",x"10",x"08",x"04",x"02",x"01",x"78",x"18",x"18",x"18",x"18",x"18",x"18",x"78",
    x"10",x"38",x"54",x"92",x"10",x"10",x"10",x"00",x"08",x"10",x"20",x"7E",x"20",x"10",x"08",x"00",
    x"08",x"04",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"7C",x"0C",x"7C",x"6C",x"7E",x"00",
    x"70",x"30",x"3E",x"36",x"36",x"36",x"3E",x"00",x"00",x"00",x"7E",x"66",x"60",x"60",x"7E",x"00",
    x"0E",x"0C",x"7C",x"6C",x"6C",x"6C",x"7C",x"00",x"00",x"00",x"7E",x"66",x"7E",x"60",x"7E",x"00",
    x"00",x"3E",x"30",x"7C",x"30",x"30",x"30",x"00",x"00",x"00",x"7E",x"6C",x"6C",x"7C",x"0C",x"7C",
    x"60",x"60",x"7C",x"6C",x"6C",x"6C",x"6E",x"00",x"18",x"00",x"38",x"18",x"18",x"18",x"7E",x"00",
    x"06",x"00",x"06",x"06",x"06",x"36",x"36",x"3E",x"60",x"60",x"66",x"6C",x"78",x"66",x"66",x"00",
    x"38",x"18",x"18",x"18",x"18",x"18",x"7E",x"00",x"00",x"00",x"FE",x"D6",x"D6",x"D6",x"D6",x"00",
    x"00",x"00",x"7E",x"36",x"36",x"36",x"36",x"00",x"00",x"00",x"7E",x"66",x"66",x"66",x"7E",x"00",
    x"00",x"00",x"7E",x"36",x"36",x"3E",x"30",x"30",x"00",x"00",x"7C",x"6C",x"6C",x"7C",x"0C",x"0E",
    x"00",x"00",x"7E",x"36",x"30",x"30",x"30",x"00",x"00",x"00",x"7E",x"60",x"7E",x"06",x"7E",x"00",
    x"00",x"30",x"7E",x"30",x"30",x"30",x"3E",x"00",x"00",x"00",x"6C",x"6C",x"6C",x"6C",x"7E",x"00",
    x"00",x"00",x"66",x"66",x"66",x"3C",x"18",x"00",x"00",x"00",x"D6",x"D6",x"D6",x"FE",x"6C",x"00",
    x"00",x"00",x"66",x"3C",x"18",x"3C",x"66",x"00",x"00",x"00",x"76",x"36",x"36",x"3E",x"06",x"3E",
    x"00",x"00",x"7E",x"06",x"18",x"60",x"7E",x"00",x"0E",x"08",x"08",x"30",x"08",x"08",x"0E",x"00",
    x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"70",x"10",x"10",x"0C",x"10",x"10",x"70",x"00",
    x"00",x"00",x"00",x"78",x"1E",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"00",x"00",x"00",x"00",x"00",x"03",x"1F",x"FF",x"00",x"00",x"00",x"00",x"00",x"C0",x"F8",x"FF",
    x"FF",x"1F",x"03",x"00",x"00",x"00",x"00",x"00",x"FF",x"F8",x"C0",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"01",x"0F",x"7F",x"FF",x"FF",x"FF",x"00",x"00",x"80",x"F0",x"FE",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"7F",x"0F",x"01",x"00",x"00",x"FF",x"FF",x"FF",x"FE",x"F0",x"80",x"00",x"00",
    x"07",x"3F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E0",x"FC",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"3F",x"07",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FC",x"E0",
    x"00",x"00",x"00",x"00",x"03",x"0F",x"3F",x"FF",x"00",x"00",x"00",x"00",x"C0",x"F0",x"FC",x"FF",
    x"FF",x"3F",x"0F",x"03",x"00",x"00",x"00",x"00",x"FF",x"FC",x"F0",x"C0",x"00",x"00",x"00",x"00",
    x"03",x"0F",x"3F",x"FF",x"FF",x"FF",x"FF",x"FF",x"C0",x"F0",x"FC",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"3F",x"0F",x"03",x"FF",x"FF",x"FF",x"FF",x"FF",x"FC",x"F0",x"C0",
    x"01",x"03",x"07",x"0F",x"1F",x"3F",x"7F",x"FF",x"80",x"C0",x"E0",x"F0",x"F8",x"FC",x"FE",x"FF",
    x"FF",x"7F",x"3F",x"1F",x"0F",x"07",x"03",x"01",x"FF",x"FE",x"FC",x"F8",x"F0",x"E0",x"C0",x"80",
    x"00",x"00",x"00",x"00",x"01",x"03",x"07",x"0F",x"00",x"00",x"00",x"00",x"80",x"C0",x"E0",x"F0",
    x"0F",x"07",x"03",x"01",x"00",x"00",x"00",x"00",x"F0",x"E0",x"C0",x"80",x"00",x"00",x"00",x"00",
    x"1F",x"3F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FF",x"F8",x"FC",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"7F",x"3F",x"1F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FC",x"F8",
    x"1F",x"1F",x"3F",x"3F",x"7F",x"7F",x"FF",x"FF",x"F8",x"F8",x"FC",x"FC",x"FE",x"FE",x"FF",x"FF",
    x"FF",x"FF",x"7F",x"7F",x"3F",x"3F",x"1F",x"1F",x"FF",x"FF",x"FE",x"FE",x"FC",x"FC",x"F8",x"F8",
    x"01",x"01",x"03",x"03",x"07",x"07",x"0F",x"0F",x"80",x"80",x"C0",x"C0",x"E0",x"E0",x"F0",x"F0",
    x"0F",x"0F",x"07",x"07",x"03",x"03",x"01",x"01",x"F0",x"F0",x"E0",x"E0",x"C0",x"C0",x"80",x"80",
    x"3F",x"3F",x"7F",x"7F",x"7F",x"FF",x"FF",x"FF",x"FC",x"FC",x"FE",x"FE",x"FE",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"7F",x"7F",x"7F",x"3F",x"3F",x"FF",x"FF",x"FF",x"FE",x"FE",x"FE",x"FC",x"FC",
    x"07",x"0F",x"0F",x"0F",x"1F",x"1F",x"1F",x"3F",x"E0",x"F0",x"F0",x"F0",x"F8",x"F8",x"F8",x"FC",
    x"3F",x"1F",x"1F",x"1F",x"0F",x"0F",x"0F",x"07",x"FC",x"F8",x"F8",x"F8",x"F0",x"F0",x"F0",x"E0",
    x"01",x"01",x"01",x"03",x"03",x"03",x"07",x"07",x"80",x"80",x"80",x"C0",x"C0",x"C0",x"E0",x"E0",
    x"07",x"07",x"03",x"03",x"03",x"01",x"01",x"01",x"E0",x"E0",x"C0",x"C0",x"C0",x"80",x"80",x"80",
    x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"FF",
    x"00",x"00",x"00",x"00",x"0F",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"F0",x"FF",x"FF",x"FF",
    x"00",x"00",x"0F",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"F0",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"0F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"01",x"01",x"01",x"01",x"03",x"03",x"03",x"03",x"80",x"80",x"80",x"80",x"C0",x"C0",x"C0",x"C0",
    x"07",x"07",x"07",x"07",x"0F",x"0F",x"0F",x"0F",x"E0",x"E0",x"E0",x"E0",x"F0",x"F0",x"F0",x"F0",
    x"1F",x"1F",x"1F",x"1F",x"3F",x"3F",x"3F",x"3F",x"F8",x"F8",x"F8",x"F8",x"FC",x"FC",x"FC",x"FC",
    x"7F",x"7F",x"7F",x"7F",x"FF",x"FF",x"FF",x"FF",x"FE",x"FE",x"FE",x"FE",x"FF",x"FF",x"FF",x"FF",
    x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"0F",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0",
    x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"F0",x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"0F",
    x"00",x"00",x"00",x"00",x"0F",x"F0",x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"0F",x"00",x"00",
    x"00",x"00",x"0F",x"F0",x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"0F",x"00",x"00",x"00",x"00",
    x"0F",x"F0",x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"03",x"1C",x"E0",x"00",x"00",x"00",x"00",x"00",x"C0",x"38",x"07",
    x"00",x"00",x"01",x"0E",x"70",x"80",x"00",x"00",x"00",x"00",x"80",x"70",x"0E",x"01",x"00",x"00",
    x"07",x"38",x"C0",x"00",x"00",x"00",x"00",x"00",x"E0",x"1C",x"03",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"03",x"0C",x"30",x"C0",x"00",x"00",x"00",x"00",x"C0",x"30",x"0C",x"03",
    x"03",x"0C",x"30",x"C0",x"00",x"00",x"00",x"00",x"C0",x"30",x"0C",x"03",x"00",x"00",x"00",x"00",
    x"10",x"20",x"40",x"80",x"00",x"00",x"00",x"00",x"08",x"04",x"02",x"01",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"80",x"40",x"20",x"10",x"00",x"00",x"00",x"00",x"01",x"02",x"04",x"08",
    x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
    x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",x"0C",
    x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",
    x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"08",x"08",x"08",x"08",x"08",x"08",x"08",x"08",
    x"F0",x"F0",x"F0",x"F0",x"00",x"00",x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"F0",x"F0",x"F0",x"F0",x"00",x"00",x"00",x"00",x"0F",x"0F",x"0F",x"0F",
    x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",
    x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
    x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"7E",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",
    x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"4D",x"61",x"74",x"74",x"65",x"6C",x"20",x"45",
    x"6C",x"65",x"63",x"74",x"72",x"6F",x"6E",x"69",x"63",x"73",x"20",x"20",x"20",x"20",x"20",x"20",
    x"20",x"70",x"72",x"65",x"73",x"65",x"6E",x"74",x"73",x"00",x"43",x"6F",x"70",x"72",x"20",x"40",
    x"20",x"31",x"39",x"38",x"34",x"20",x"4D",x"61",x"74",x"74",x"65",x"6C",x"00",x"FF",x"FF",x"24",
    x"00",x"82",x"AE",x"08",x"C9",x"10",x"14",x"88",x"91",x"08",x"42",x"22",x"02",x"82",x"18",x"89",
    x"08",x"20",x"8A",x"23",x"02",x"02",x"20",x"B8",x"82",x"28",x"0A",x"20",x"AE",x"20",x"8A",x"AA",
    x"92",x"20",x"8A",x"B8",x"82",x"88",x"22",x"B8",x"82",x"88",x"EA",x"8A",x"AA",x"AE",x"88",x"68",
    x"AE",x"0C",x"27",x"11",x"1F",x"00",x"2B",x"32",x"0A",x"4A",x"D1",x"B8",x"04",x"51",x"72",x"6A",
    x"10",x"2C",x"05",x"42",x"62",x"62",x"7C",x"F0",x"2C",x"0E",x"00",x"34",x"04",x"00",x"C3",x"98",
    x"B8",x"04",x"C0",x"C3",x"42",x"4D",x"D1",x"C0",x"14",x"60",x"0C",x"02",x"B8",x"00",x"04",x"00",
    x"DC",x"59",x"29",x"0A",x"59",x"09",x"08",x"04",x"00",x"DC",x"59",x"29",x"05",x"20",x"15",x"14",
    x"60",x"0C",x"05",x"89",x"04",x"0A",x"B8",x"00",x"04",x"00",x"DC",x"59",x"29",x"0E",x"20",x"26",
    x"4F",x"43",x"5F",x"0A",x"1A",x"BC",x"E8",x"A5",x"A1",x"B9",x"FF",x"04",x"0D",x"B8",x"08",x"10",
    x"71",x"29",x"03",x"71",x"0F",x"69",x"10",x"23",x"03",x"41",x"69",x"7D",x"F0",x"2C",x"16",x"5B",
    x"09",x"10",x"BC",x"E8",x"A5",x"A1",x"B8",x"04",x"7D",x"56",x"10",x"2C",x"04",x"6A",x"7D",x"F0",
    x"2C",x"0C",x"5B",x"09",x"0D",x"BC",x"E8",x"A5",x"BA",x"EF",x"A0",x"91",x"69",x"50",x"12",x"62",
    x"2E",x"07",x"5B",x"09",x"0A",x"BC",x"E8",x"A5",x"A1",x"19",x"69",x"7D",x"F0",x"2C",x"06",x"5B",
    x"09",x"1A",x"B8",x"08",x"BC",x"E8",x"A5",x"A1",x"79",x"72",x"69",x"7D",x"F0",x"2C",x"07",x"42",
    x"72",x"10",x"2C",x"0F",x"BC",x"E8",x"B1",x"61",x"7C",x"F0",x"2C",x"05",x"B3",x"BC",x"E8",x"B5",
    x"A0",x"68",x"7C",x"F0",x"2C",x"05",x"B0",x"10",x"0C",x"01",x"B5",x"B7",x"C0",x"60",x"7C",x"F0",
    x"2C",x"04",x"3C",x"08",x"8B",x"BB",x"00",x"04",x"03",x"D9",x"4B",x"D9",x"8B",x"BB",x"C0",x"D9",
    x"4F",x"43",x"7A",x"53",x"AF",x"7C",x"F0",x"24",x"98",x"75",x"85",x"E5",x"14",x"65",x"B7",x"00");

  CONSTANT INIT_ECS : arr16 := (
    x"02BA",x"017F",x"0001",x"02BB",x"000F",x"0070",x"0004",x"0120",
    x"001F",x"037A",x"0170",x"020C",x"0003",x"0004",x"0370",x"0026",
    x"02A0",x"0150",x"020C",x"0007",x"03BA",x"00F0",x"0001",x"033C",
    x"0000",x"0010",x"00A7",x"0013",x"0012",x"0220",x"0018",x"009C",
    x"02B9",x"0294",x"004D",x"01E1",x"00A0",x"03B8",x"000F",x"0001",
    x"03F8",x"00FF",x"000F",x"01C4",x"0261",x"0014",x"00AF",x"0275",
    x"0281",x"02F0",x"0339",x"0008",x"0288",x"0080",x"020B",x"0002",
    x"03B8",x"0200",x"02B7",x"0275",x"0004",x"0174",x"01F2",x"0001",
    x"02BC",x"00B1",x"0040",x"02A2",x"00E2",x"033A",x"0003",x"02B8",
    x"000D",x"0250",x"02B8",x"0010",x"0004",x"01EC",x"03E0",x"02A0",
    x"0081",x"03B8",x"00E0",x"0378",x"00A0",x"020C",x"0018",x"03B9",
    x"001F",x"0009",x"00F9",x"02CF",x"0080",x"010E",x"007D",x"007D",
    x"007D",x"0195",x"01C9",x"010B",x"0160",x"0131",x"007A",x"025C",
    x"017C",x"029F",x"0278",x"0281",x"026D",x"0030",x"0195",x"0004",
    x"0120",x"03C9",x"0004",x"01EC",x"0049",x"02B9",x"0082",x"02A0",
    x"0141",x"0204",x"0006",x"02A0",x"0148",x"0204",x"0002",x"02FC",
    x"0005",x"0004",x"0120",x"031A",x"0004",x"0174",x"01D4",x"0004",
    x"0178",x"00AF",x"0200",x"004D",x"02A0",x"0378",x"000D",x"0204",
    x"0048",x"0001",x"02BD",x"00E9",x"0047",x"0001",x"02A9",x"0089",
    x"020C",x"000A",x"0001",x"02B9",x"00FE",x"0025",x"0004",x"0120",
    x"0399",x"000C",x"0220",x"0017",x"0274",x"0271",x"02AA",x"0093",
    x"004A",x"00D3",x"004A",x"00D3",x"00D9",x"02F9",x"0003",x"0004",
    x"0120",x"0399",x"02B1",x"0011",x"0288",x"02FB",x"0012",x"0158",
    x"0203",x"0013",x"0009",x"008C",x"0004",x"0174",x"028B",x"0080",
    x"020C",x"0004",x"01E4",x"0004",x"0174",x"028B",x"0004",x"0174",
    x"0292",x"02B4",x"000C",x"0220",x"0040",x"0001",x"02B9",x"00EB",
    x"0047",x"0288",x"0008",x"0248",x"0220",x"000C",x"0004",x"0174",
    x"01B3",x"02B8",x"0001",x"02B7",x"0001",x"02BD",x"00B5",x"0047",
    x"0001",x"02AB",x"0013",x"0299",x"0339",x"0008",x"00CB",x"0298",
    x"0080",x"020C",x"0040",x"00A2",x"000A",x"033C",x"0002",x"00CC",
    x"0290",x"0378",x"0080",x"020C",x"0002",x"02FA",x"0005",x"000A",
    x"0290",x"0378",x"0080",x"020C",x"0004",x"02FA",x"0002",x"0200",
    x"0003",x"0004",x"0178",x"008B",x"0091",x"00A2",x"0004",x"01EC",
    x"0058",x"009A",x"0004",x"01EC",x"0058",x"02FC",x"0002",x"0001",
    x"02BA",x"00B3",x"0040",x"0272",x"0004",x"0178",x"008B",x"0094",
    x"02B2",x"000A",x"0290",x"0378",x"0080",x"020C",x"0004",x"02FA",
    x"0002",x"0200",x"0003",x"0004",x"0178",x"008B",x"0091",x"00A2",
    x"0004",x"01EC",x"0058",x"0001",x"02BD",x"00B1",x"0040",x"02A8",
    x"0338",x"0003",x"00AA",x"000A",x"00C5",x"033D",x"0006",x"00AB",
    x"0004",x"0178",x"008B",x"0004",x"01E0",x"0308",x"0020",x"0223",
    x"0067",x"0001",x"02BD",x"00B1",x"0040",x"02A8",x"0338",x"0005",
    x"00C5",x"0001",x"02AC",x"0004",x"01EC",x"039F",x"0080",x"022B",
    x"0005",x"0204",x"0014",x"01C0",x"0200",x"0001",x"0275",x"00A1",
    x"0001",x"02BD",x"00B5",x"0047",x"0269",x"0041",x"0269",x"0080",
    x"020C",x"0004",x"0004",x"0174",x"0204",x"01C0",x"02B7",x"01C0",
    x"0010",x"02B7",x"0004",x"01EC",x"0049",x"02B8",x"0001",x"0283",
    x"035C",x"0004",x"01EC",x"0340",x"00A2",x"0272",x"0004",x"0178",
    x"008B",x"0272",x"0093",x"01C0",x"0004",x"01E0",x"0059",x"02B2",
    x"0281",x"035C",x"0004",x"01EC",x"0058",x"02B3",x"000B",x"009D",
    x"0001",x"02A9",x"01C0",x"0220",x"0034",x"0281",x"015D",x"03B9",
    x"0004",x"0204",x"0008",x"0001",x"02BD",x"00B5",x"0047",x"0001",
    x"02AB",x"0200",x"0001",x"01DB",x"0001",x"02B9",x"00C2",x"0047",
    x"028A",x"037A",x"0005",x"020B",x"000B",x"009D",x"033D",x"0003",
    x"0001",x"02AB",x"009A",x"0004",x"012C",x"01DE",x"0220",x"00D6",
    x"004A",x"0001",x"02FA",x"00B8",x"0047",x"0253",x"000A",x"0043",
    x"0253",x"028A",x"000A",x"024A",x"00A5",x"0001",x"02AA",x"01E4",
    x"0004",x"01EC",x"039F",x"0142",x"0204",x"0004",x"0080",x"022C",
    x"0008",x"02B7",x"0281",x"015D",x"03B9",x"0004",x"020C",x"0005",
    x"0274",x"0004",x"0174",x"0212",x"02B4",x"01C0",x"0220",x"0080",
    x"0001",x"02B9",x"00C2",x"0047",x"028A",x"0092",x"0224",x"0078",
    x"0012",x"024A",x"004A",x"0001",x"02FA",x"00B8",x"0047",x"0095",
    x"0001",x"02AC",x"00A4",x"0224",x"0085",x"02B8",x"0001",x"0220",
    x"0099",x"0004",x"0174",x"03F9",x"02A0",x"0270",x"0091",x"0001",
    x"02BA",x"00C6",x"0047",x"0272",x"0004",x"01EC",x"0058",x"0004",
    x"0174",x"03F9",x"02B3",x"0274",x"0004",x"01E0",x"0308",x"0020",
    x"02B5",x"02B1",x"03B9",x"0003",x"0339",x"0002",x"0148",x"022C",
    x"0137",x"0284",x"0354",x"02FC",x"002C",x"02A2",x"00A3",x"00E2",
    x"033A",x"0002",x"02A8",x"0260",x"016A",x"022C",x"0004",x"01C0",
    x"0268",x"009C",x"0012",x"0220",x"01DA",x"0004",x"0120",x"03C9",
    x"0004",x"0120",x"0380",x"02A0",x"0378",x"000D",x"0224",x"0156",
    x"0274",x"0283",x"0354",x"009D",x"01C0",x"0268",x"0001",x"037D",
    x"0099",x"0040",x"022C",x"0006",x"02B4",x"0273",x"0014",x"0004",
    x"0120",x"031A",x"02B3",x"0001",x"02BA",x"00B7",x"0047",x"0292",
    x"03BA",x"0010",x"0204",x"0018",x"0274",x"009C",x"01C0",x"02B9",
    x"0001",x"02BA",x"0002",x"0283",x"035C",x"029D",x"03BD",x"0080",
    x"020C",x"0003",x"02BB",x"0020",x"0263",x"0004",x"0120",x"03EE",
    x"00A3",x"02B4",x"0200",x"002B",x"0274",x"0273",x"0004",x"0124",
    x"019D",x"0001",x"02BA",x"00B7",x"0047",x"0292",x"0091",x"03BA",
    x"0007",x"0093",x"0080",x"0203",x"0001",x"01C0",x"00C3",x"02FB",
    x"0003",x"03B9",x"0008",x"02BD",x"0009",x"0089",x"0204",x"0002",
    x"02FD",x"000A",x"015D",x"0203",x"0004",x"02B3",x"02B4",x"0220",
    x"003C",x"011D",x"02B4",x"00EC",x"01C9",x"0220",x"003B",x"0001",
    x"02B9",x"00B7",x"0047",x"0289",x"03B9",x"0008",x"0204",x"000B",
    x"000C",x"0274",x"02B8",x"000D",x"0258",x"0004",x"012C",x"02DE",
    x"02B4",x"0220",x"0077",x"000C",x"0001",x"037B",x"0090",x"0040",
    x"0223",x"0010",x"02A0",x"0378",x"000D",x"020C",x"0003",x"0014",
    x"0220",x"0018",x"0001",x"02BB",x"008F",x"0040",x"0220",x"007A",
    x"0004",x"0120",x"0380",x"02A0",x"0378",x"000D",x"0224",x"01E6",
    x"0001",x"033C",x"00AF",x"0040",x"0001",x"02B9",x"00FA",x"0047",
    x"024C",x"0280",x"015D",x"03B8",x"00E7",x"03F8",x"0018",x"0240",
    x"015D",x"02B5",x"02B5",x"02B7",x"02A1",x"0004",x"0120",x"03A3",
    x"0004",x"0120",x"03AE",x"0220",x"0203",x"02A1",x"0004",x"0120",
    x"03A3",x"008C",x"0281",x"0354",x"0004",x"0120",x"03AE",x"02B8",
    x"000D",x"0260",x"0001",x"02B9",x"0098",x"0040",x"0288",x"0378",
    x"0020",x"020C",x"0003",x"02B8",x"000D",x"0248",x"0004",x"012C",
    x"02DE",x"0220",x"0221",x"02BA",x"000C",x"02B8",x"000A",x"0004",
    x"01EC",x"03E0",x"02A1",x"014A",x"020B",x"0007",x"0001",x"02BC",
    x"0019",x"0027",x"0011",x"0200",x"0008",x"0011",x"0111",x"0285",
    x"02F0",x"02FD",x"000E",x"0001",x"02AC",x"0049",x"00CC",x"0001",
    x"02A1",x"008F",x"0275",x"0004",x"01EC",x"0049",x"0004",x"0174",
    x"03DF",x"0080",x"020C",x"000B",x"0004",x"0174",x"03F9",x"0091",
    x"0282",x"035C",x"0004",x"01EC",x"0058",x"0200",x"0050",x"0274",
    x"0004",x"0174",x"034B",x"0080",x"0203",x"0021",x"0008",x"0203",
    x"000B",x"0004",x"0174",x"03F9",x"0091",x"0282",x"035C",x"02FA",
    x"0015",x"0004",x"01EC",x"0058",x"0284",x"035C",x"00A5",x"02FD",
    x"0015",x"00AA",x"02BB",x"0007",x"02A0",x"02A9",x"0014",x"0015",
    x"0261",x"0268",x"0013",x"022C",x"0008",x"0200",x"001A",x"0080",
    x"0204",x"0014",x"0281",x"035C",x"008A",x"02FA",x"0015",x"0004",
    x"01EC",x"005C",x"0004",x"01EC",x"0049",x"0004",x"0174",x"03F9",
    x"0091",x"0282",x"035C",x"0004",x"01EC",x"0058",x"0004",x"0174",
    x"03F9",x"0093",x"02B4",x"02A2",x"0274",x"0004",x"0178",x"0095",
    x"02B4",x"0004",x"0174",x"03DF",x"0080",x"022C",x"004F",x"02B7",
    x"0275",x"0285",x"0354",x"02A0",x"0378",x"0001",x"0204",x"0003",
    x"0268",x"0220",x"0007",x"0280",x"0354",x"0145",x"0204",x"0008",
    x"02B8",x"000D",x"0268",x"0274",x"0004",x"012C",x"02DE",x"02B4",
    x"02B7",x"0275",x"00A2",x"0012",x"0004",x"0178",x"008B",x"0004",
    x"01EC",x"0058",x"02B7",x"0275",x"0011",x"004D",x"008D",x"004D",
    x"00E9",x"0001",x"02F9",x"0075",x"0047",x"02B7",x"0275",x"008D",
    x"02F9",x"0014",x"02A0",x"0378",x"0001",x"0204",x"0008",x"0378",
    x"000D",x"0204",x"0004",x"0268",x"0169",x"022C",x"000C",x"014D",
    x"020C",x"0002",x"00AC",x"02B7",x"02B8",x"0020",x"0268",x"0220",
    x"0009",x"0275",x"000A",x"0274",x"0014",x"00A5",x"01DB",x"0162",
    x"0204",x"001A",x"02A0",x"009B",x"020C",x"0012",x"0378",x"0080",
    x"020C",x"0004",x"02BB",x"0005",x"0200",x"000B",x"0378",x"0084",
    x"0224",x"0012",x"0378",x"008A",x"0224",x"0016",x"0200",x"0001",
    x"0013",x"0268",x"0220",x"001C",x"02B4",x"02B7",x"0275",x"0285",
    x"015D",x"03BD",x"007F",x"03FD",x"0080",x"0245",x"015D",x"0270",
    x"0271",x"0272",x"0281",x"035C",x"0001",x"02BA",x"00EE",x"0047",
    x"0004",x"01EC",x"005C",x"0095",x"00A2",x"026A",x"0042",x"026A",
    x"008B",x"02B2",x"02B1",x"02B0",x"0268",x"026A",x"029D",x"03BD",
    x"0080",x"0204",x"0007",x"029D",x"03BD",x"007F",x"025D",x"02BD",
    x"002D",x"0265",x"0270",x"0271",x"0272",x"0281",x"035C",x"008A",
    x"033A",x"0007",x"0004",x"01EC",x"005C",x"02B2",x"02B1",x"02B0",
    x"0089",x"0204",x"0037",x"0270",x"0272",x"0271",x"0004",x"0124",
    x"019D",x"0083",x"02B1",x"02B2",x"02B0",x"0103",x"009D",x"009B",
    x"0203",x"0005",x"0023",x"0001",x"03FB",x"0000",x"0040",x"0379",
    x"0002",x"020C",x"0004",x"0001",x"03FB",x"0000",x"0080",x"0273",
    x"0270",x"0272",x"00A8",x"0020",x"0004",x"01EC",x"006A",x"0001",
    x"02BB",x"00C6",x"0047",x"0273",x"0004",x"01E0",x"00BB",x"02B2",
    x"0091",x"02F9",x"0007",x"0004",x"01EC",x"005C",x"02B2",x"02B0",
    x"0200",x"0003",x"02BB",x"00FF",x"0273",x"01C9",x"0011",x"0080",
    x"0203",x"0004",x"02BB",x"002E",x"0263",x"01C9",x"0001",x"02BD",
    x"00C3",x"0047",x"026A",x"0269",x"0270",x"0004",x"01EC",x"006A",
    x"0281",x"035C",x"008A",x"02FA",x"0015",x"0004",x"01EC",x"005C",
    x"008A",x"0339",x"0007",x"0004",x"01EC",x"005C",x"0093",x"0273",
    x"02FB",x"000E",x"0004",x"01E0",x"0267",x"02B3",x"033B",x"0007",
    x"0004",x"01E4",x"01A2",x"0378",x"000A",x"020B",x"0002",x"02B8",
    x"0009",x"0083",x"02FB",x"0030",x"0263",x"0080",x"0204",x"001F",
    x"0283",x"035C",x"0004",x"01EC",x"0340",x"0273",x"02FB",x"0015",
    x"0004",x"01E0",x"00BB",x"02B1",x"028A",x"03FA",x"0080",x"024A",
    x"008B",x"033B",x"0007",x"0273",x"01C0",x"0004",x"01E0",x"0059",
    x"02B2",x"0091",x"02F9",x"0007",x"0004",x"01EC",x"005C",x"02B0",
    x"0001",x"02BD",x"00C3",x"0047",x"02AA",x"02A9",x"0379",x"00FF",
    x"020C",x"0002",x"01C9",x"0011",x"0010",x"0223",x"0060",x"0089",
    x"0203",x"0009",x"01C9",x"014A",x"0204",x"0006",x"02BB",x"002E",
    x"0263",x"0200",x"0001",x"0009",x"014A",x"022C",x"0070",x"0004",
    x"01EC",x"006A",x"0001",x"02BB",x"00E2",x"0047",x"02B8",x"0005",
    x"0004",x"01EC",x"0340",x"0273",x"0004",x"01E0",x"00BB",x"02B8",
    x"0001",x"02B3",x"033B",x"001C",x"0273",x"0004",x"01E0",x"0059",
    x"02B1",x"02F9",x"0007",x"0288",x"03B8",x"0080",x"0204",x"0017",
    x"00A2",x"0012",x"0290",x"0378",x"002E",x"0224",x"0005",x"0004",
    x"012C",x"01D2",x"0201",x"004A",x"0008",x"0378",x"003A",x"020C",
    x"0005",x"02B8",x"0030",x"0250",x"0220",x"0014",x"0250",x"02B0",
    x"0378",x"00FF",x"0204",x"0033",x"02B9",x"0045",x"0261",x"0083",
    x"009D",x"0001",x"03BB",x"0000",x"0040",x"0001",x"03BD",x"0000",
    x"0080",x"009B",x"0204",x"0005",x"02B9",x"002D",x"0261",x"0200",
    x"0006",x"02B9",x"0020",x"0034",x"0034",x"0034",x"0261",x"03B8",
    x"00FF",x"0034",x"0083",x"0081",x"02BA",x"000A",x"0004",x"011C",
    x"01FB",x"0081",x"02F8",x"0030",x"0260",x"02B8",x"000A",x"0004",
    x"011C",x"01DC",x"0113",x"0098",x"02F8",x"0030",x"0260",x"02B8",
    x"0007",x"0004",x"0114",x"02DB",x"015D",x"02B7",x"02B0",x"0378",
    x"00FF",x"0204",x"0021",x"000A",x"0291",x"0379",x"002E",x"020C",
    x"0001",x"000A",x"02B9",x"0031",x"0251",x"0085",x"0040",x"03B8",
    x"0040",x"0204",x"0002",x"0015",x"0015",x"000D",x"0275",x"000A",
    x"0290",x"0378",x"002E",x"0224",x"0005",x"0004",x"012C",x"01D2",
    x"0229",x"000A",x"0220",x"0064",x"0282",x"035C",x"0001",x"02B9",
    x"00EE",x"0047",x"0004",x"01EC",x"005C",x"008D",x"02FD",x"0007",
    x"0001",x"02AC",x"02A8",x"02AA",x"0008",x"0085",x"00D5",x"0014",
    x"01C9",x"037D",x"0007",x"022B",x"01A5",x"000C",x"01C0",x"02B9",
    x"0001",x"02BA",x"0002",x"0220",x"01AD",x"0275",x"0274",x"02B8",
    x"0007",x"0004",x"0114",x"02E6",x"015D",x"0004",x"0170",x"00A2",
    x"0204",x"004C",x"0288",x"0270",x"03B8",x"007F",x"0248",x"008A",
    x"02FA",x"0015",x"0004",x"01EC",x"005C",x"0004",x"01E0",x"01DD",
    x"0090",x"008B",x"0004",x"01E4",x"01FB",x"0273",x"0001",x"02BB",
    x"0067",x"0026",x"0004",x"01E0",x"00BB",x"02B3",x"02BC",x"004B",
    x"0004",x"01E4",x"01DC",x"0270",x"0024",x"0160",x"0204",x"001B",
    x"0004",x"01EC",x"006A",x"0281",x"035C",x"0288",x"03F8",x"0080",
    x"0248",x"01C0",x"008B",x"0273",x"02FB",x"0015",x"0004",x"01E0",
    x"0059",x"02B1",x"0288",x"03B8",x"0080",x"0204",x"0004",x"02B0",
    x"0010",x"0220",x"001F",x"008A",x"02F9",x"0015",x"0004",x"01EC",
    x"005C",x"02B0",x"02B1",x"033A",x"0007",x"0251",x"0285",x"015D",
    x"03BD",x"007F",x"0245",x"015D",x"02B4",x"02B7",x"0040",x"0000",
    x"0000",x"0000",x"0000",x"0000",x"0000",x"0041",x"00A0",x"0000",
    x"0000",x"0000",x"0000",x"0000",x"0042",x"0064",x"0000",x"0000",
    x"0000",x"0000",x"0000",x"0044",x"0027",x"0010",x"0000",x"0000",
    x"0000",x"0000",x"0047",x"005F",x"005E",x"0010",x"0000",x"0000",
    x"0000",x"004E",x"0023",x"0086",x"00F2",x"006F",x"00C1",x"0000",
    x"005B",x"004E",x"00E2",x"00D6",x"00D4",x"0015",x"00B8",x"0076",
    x"0018",x"004F",x"0003",x"00E9",x"003F",x"00FA",x"0040",x"0019",
    x"0099",x"0099",x"0099",x"0099",x"009A",x"0001",x"0028",x"00F5",
    x"00C2",x"008F",x"005C",x"0029",x"0003",x"0068",x"00DB",x"008B",
    x"00AC",x"0071",x"000D",x"0006",x"002A",x"00F3",x"001D",x"00C4",
    x"0061",x"0018",x"000D",x"0073",x"004A",x"00CA",x"005F",x"0062",
    x"0027",x"001A",x"0033",x"00EC",x"0047",x"00AB",x"0051",x"004E",
    x"0035",x"00A8",x"007F",x"00EA",x"0027",x"00A5",x"003A",x"0041",
    x"0013",x"0042",x"00F7",x"00F9",x"0000",x"0000",x"00FD",x"00E4",
    x"0003",x"00E5",x"000F",x"00E6",x"0016",x"00E6",x"003F",x"00E6",
    x"006C",x"00E6",x"0076",x"00E6",x"00AB",x"00E6",x"00A3",x"00E6",
    x"00AF",x"00E6",x"0035",x"00E5",x"00C2",x"00E6",x"00C2",x"00E6",
    x"00C2",x"00E6",x"00A7",x"00E6",x"005F",x"00E7",x"0043",x"00E7",
    x"0007",x"00E7",x"00FA",x"00E6",x"00D3",x"00E4",x"00D3",x"00E4",
    x"00D3",x"00E4",x"004C",x"0049",x"0053",x"0054",x"0043",x"004C",
    x"004F",x"0044",x"0043",x"0053",x"0041",x"0056",x"0044",x"0045",
    x"004C",x"0020",x"0052",x"0055",x"004E",x"0020",x"004E",x"0045",
    x"0057",x"0020",x"0043",x"0056",x"0052",x"0046",x"004D",x"0045",
    x"004E",x"0055",x"0000",x"0054",x"004F",x"004E",x"0045",x"0045",
    x"004E",x"0056",x"0054",x"004E",x"004F",x"0049",x"0053",x"0045",
    x"004E",x"0056",x"004E",x"0044",x"0049",x"0053",x"0054",x"0048",
    x"0055",x"0053",x"0048",x"004E",x"004F",x"0054",x"0045",x"0053",
    x"0048",x"004F",x"0057",x"0047",x"0052",x"0041",x"0042",x"004F",
    x"0055",x"0054",x"0050",x"004C",x"0049",x"004E",x"004B",x"0048",
    x"0041",x"004E",x"0044",x"0000",x"0058",x"0056",x"0059",x"0056",
    x"0058",x"0050",x"0059",x"0050",x"0043",x"004F",x"0052",x"004E",
    x"0056",x"0053",x"0059",x"004D",x"0058",x"0053",x"0058",x"004D",
    x"0046",x"004D",x"0041",x"0041",x"0041",x"0042",x"0041",x"0043",
    x"0059",x"0053",x"0053",x"0051",x"0050",x"0043",x"0042",x"004B",
    x"0049",x"0054",x"0041",x"0024",x"0042",x"0024",x"0043",x"0024",
    x"0000",x"002B",x"00E3",x"0041",x"00E3",x"0039",x"00E3",x"004F",
    x"00E3",x"0083",x"00E3",x"00AE",x"00E3",x"00BE",x"00E4",x"005E",
    x"00E4",x"008E",x"00E4",x"0031",x"0027",x"0047",x"00E4",x"0057",
    x"00E3",x"0001",x"02BD",x"0019",x"0047",x"02A8",x"03B8",x"0080",
    x"0281",x"015E",x"03B9",x"007F",x"01C8",x"0240",x"015E",x"02B7",
    x"0275",x"0284",x"0354",x"00A3",x"02FB",x"002A",x"0004",x"0128",
    x"021A",x"000B",x"0092",x"020C",x"000B",x"02B9",x"0010",x"0004",
    x"0128",x"0226",x"0204",x"0008",x"02F9",x"0004",x"0200",x"0004",
    x"01C9",x"0004",x"0128",x"0226",x"0089",x"0204",x"001B",x"0011",
    x"0088",x"03F8",x"00A0",x"0258",x"000B",x"0009",x"00F9",x"02CF",
    x"01C6",x"01E2",x"002F",x"003F",x"00DE",x"01F1",x"01AD",x"0262",
    x"01E9",x"01E9",x"0262",x"0180",x"0262",x"0090",x"007E",x"0079",
    x"0079",x"0184",x"0004",x"0128",x"03A0",x"0004",x"0178",x"032C",
    x"0004",x"0128",x"0293",x"02B8",x"0082",x"0004",x"0128",x"01A8",
    x"02B8",x"0082",x"0258",x"000B",x"0004",x"0178",x"01BE",x"0080",
    x"020B",x"022D",x"0004",x"0178",x"00F8",x"0200",x"0233",x"02A0",
    x"0378",x"000D",x"0204",x"022E",x"0258",x"000B",x"0001",x"02B8",
    x"0016",x"0006",x"0004",x"017C",x"039A",x"0220",x"000F",x"01D2",
    x"037A",x"0007",x"0204",x"021E",x"0004",x"012C",x"03B7",x"0378",
    x"000D",x"020C",x"0005",x"0092",x"0204",x"0209",x"0200",x"0212",
    x"0378",x"002E",x"0204",x"0009",x"0378",x"002D",x"0204",x"0005",
    x"0004",x"012C",x"01D2",x"0221",x"001C",x"0014",x"000A",x"0272",
    x"0004",x"01E8",x"02F0",x"02B2",x"02B8",x"000D",x"0258",x"000B",
    x"0004",x"012C",x"03B7",x"0378",x"000D",x"0204",x"01F3",x"0378",
    x"002C",x"022C",x"000A",x"0014",x"0004",x"0128",x"01A8",x"0220",
    x"0038",x"0004",x"012C",x"0024",x"0200",x"01E4",x"0004",x"012C",
    x"0024",x"0004",x"0128",x"03A0",x"02B8",x"0082",x"0004",x"0128",
    x"01A8",x"02BA",x"0014",x"0004",x"0128",x"03DE",x"0200",x"01D2",
    x"0004",x"012C",x"03B7",x"0014",x"02BA",x"000C",x"02B8",x"0002",
    x"0004",x"01EC",x"03E0",x"0272",x"0004",x"0120",x"002F",x"0204",
    x"000F",x"020B",x"000D",x"008D",x"02FD",x"0014",x"0001",x"02A9",
    x"02BA",x"0004",x"0004",x"0128",x"0264",x"0089",x"020C",x"000E",
    x"0001",x"02B9",x"00BB",x"0026",x"02BA",x"0004",x"0004",x"0128",
    x"0264",x"0089",x"0204",x"019A",x"0200",x"001A",x"0011",x"0065",
    x"02B2",x"00D1",x"0009",x"0259",x"000B",x"01D2",x"033C",x"0003",
    x"0001",x"02B8",x"0002",x"0007",x"0004",x"017C",x"039A",x"000A",
    x"000C",x"037A",x"0004",x"022C",x"0008",x"0014",x"0200",x"018A",
    x"0011",x"0065",x"02B5",x"0220",x"001A",x"0034",x"0004",x"0128",
    x"03A0",x"0004",x"0178",x"032C",x"0001",x"02BC",x"0087",x"0040",
    x"02A0",x"0378",x"000D",x"0204",x"016A",x"0378",x"00CB",x"022B",
    x"0008",x"0378",x"00CE",x"0223",x"000C",x"0014",x"0274",x"0273",
    x"02A2",x"0285",x"0354",x"02FD",x"002A",x"0001",x"02AB",x"01E4",
    x"0004",x"01EC",x"039F",x"0204",x"0063",x"022B",x"0006",x"00A5",
    x"02A9",x"0379",x"00A4",x"022C",x"000C",x"02A9",x"014A",x"022C",
    x"0010",x"0143",x"0204",x"0004",x"02B3",x"02B4",x"0200",x"013F",
    x"0004",x"012C",x"0298",x"02B3",x"02B4",x"0004",x"0128",x"02B2",
    x"01C0",x"0001",x"02BB",x"00B4",x"0040",x"0273",x"0299",x"0379",
    x"0080",x"020C",x"0005",x"02FB",x"0002",x"0004",x"01E4",x"01A2",
    x"0378",x"0001",x"0203",x"0002",x"02B8",x"0001",x"0378",x"00FB",
    x"020B",x"0002",x"02B8",x"00FA",x"0081",x"004D",x"0001",x"02BD",
    x"0007",x"0041",x"0001",x"02AA",x"0001",x"02AB",x"0094",x"00CC",
    x"02FC",x"0005",x"0163",x"0203",x"0003",x"02B3",x"0200",x"0107",
    x"0282",x"0354",x"02FA",x"002E",x"0292",x"03BA",x"001F",x"033A",
    x"000B",x"010B",x"0001",x"02BD",x"0004",x"0041",x"00D5",x"0065",
    x"0269",x"009A",x"0004",x"012C",x"03BE",x"02B3",x"0200",x"00FA",
    x"0001",x"02FA",x"0039",x"0040",x"0293",x"01C0",x"0250",x"009A",
    x"004E",x"0001",x"02BD",x"0009",x"0041",x"0001",x"02A8",x"00D0",
    x"033D",x"0002",x"0268",x"0040",x"0268",x"0220",x"0063",x"0034",
    x"01D2",x"0004",x"0128",x"03DE",x"02A0",x"0378",x"000D",x"0204",
    x"00D9",x"0014",x"0004",x"0128",x"03A0",x"02A0",x"0378",x"000D",
    x"020C",x"0003",x"0004",x"0128",x"010B",x"0378",x"0041",x"022B",
    x"000B",x"0378",x"005B",x"0223",x"000F",x"0014",x"0004",x"0128",
    x"01B6",x"0220",x"0015",x"02B8",x"000D",x"0258",x"000B",x"02A1",
    x"0089",x"0204",x"00B7",x"0088",x"00AF",x"01D2",x"0004",x"0128",
    x"03DE",x"0004",x"0128",x"03A0",x"0004",x"0178",x"032C",x"0004",
    x"0178",x"01BE",x"0080",x"020B",x"00A5",x"0004",x"0178",x"00F8",
    x"0004",x"0128",x"010B",x"0014",x"0220",x"0011",x"0004",x"0128",
    x"01B6",x"02B8",x"003D",x"0004",x"0128",x"01A8",x"0004",x"0128",
    x"01F2",x"02B8",x"0054",x"0004",x"0128",x"01A8",x"02B8",x"004F",
    x"0004",x"0128",x"01A8",x"0004",x"0128",x"01F2",x"02FB",x"0006",
    x"0200",x"0080",x"0004",x"0128",x"01B6",x"02FB",x"0002",x"0200",
    x"0079",x"0004",x"0128",x"021A",x"0092",x"0204",x"0068",x"0200",
    x"0071",x"0004",x"0128",x"03A0",x"0004",x"0178",x"032C",x"02B8",
    x"0084",x"0004",x"0128",x"01A8",x"0004",x"012C",x"004B",x"02A1",
    x"0379",x"000D",x"0204",x"0053",x"0379",x"0081",x"022B",x"0008",
    x"0379",x"0084",x"0223",x"000C",x"0259",x"000B",x"02B8",x"0006",
    x"0004",x"017C",x"039A",x"0004",x"012C",x"004B",x"02B8",x"008A",
    x"0004",x"0128",x"01A8",x"02B9",x"0018",x"0004",x"0128",x"0226",
    x"0224",x"022D",x"0001",x"02BD",x"00B2",x"0040",x"02B8",x"00B2",
    x"02F9",x"0006",x"0379",x"0013",x"0204",x"0029",x"0379",x"0009",
    x"0204",x"0004",x"0379",x"000A",x"022C",x"0241",x"0268",x"0220",
    x"0244",x"0080",x"020B",x"0003",x"0004",x"0120",x"003B",x"02B7",
    x"0275",x"02A1",x"0379",x"000D",x"0204",x"0010",x"0148",x"022C",
    x"0007",x"02B8",x"0126",x"0004",x"037C",x"039B",x"0275",x"0274",
    x"02A1",x"0379",x"000D",x"020C",x"0023",x"02B4",x"02B5",x"0281",
    x"0354",x"02F9",x"002B",x"0288",x"03F8",x"0080",x"0248",x"0004",
    x"0128",x"0322",x"009D",x"0282",x"0354",x"02FA",x"002A",x"0091",
    x"02F9",x"0002",x"0115",x"024D",x"0095",x"0001",x"02A8",x"0081",
    x"0049",x"0061",x"0224",x"003A",x"0004",x"01E0",x"0000",x"02B7",
    x"0379",x"0041",x"022B",x"002B",x"0379",x"005B",x"0223",x"002F",
    x"0259",x"000B",x"02B8",x"0024",x"02B5",x"0004",x"017C",x"039A",
    x"01C0",x"02B7",x"0275",x"02A1",x"0379",x"000D",x"0224",x"0039",
    x"0379",x"002E",x"0204",x"000C",x"0379",x"002D",x"0204",x"0008",
    x"0270",x"0088",x"0004",x"012C",x"01D2",x"02B0",x"0201",x"0005",
    x"0014",x"0004",x"01E8",x"02F0",x"02B7",x"0379",x"0041",x"022B",
    x"001D",x"0379",x"005B",x"0223",x"0021",x"0014",x"0004",x"0128",
    x"01B6",x"02B7",x"0275",x"0273",x"0004",x"012C",x"01AE",x"02B3",
    x"025A",x"000B",x"0042",x"025A",x"000B",x"02B7",x"0275",x"02B8",
    x"000E",x"0004",x"01EC",x"03E0",x"0273",x"0001",x"02F9",x"0049",
    x"002B",x"0004",x"012C",x"03B7",x"02BA",x"0004",x"0274",x"0014",
    x"0271",x"0004",x"0128",x"0264",x"0089",x"0204",x"0021",x"02B5",
    x"02B4",x"0015",x"008B",x"00EB",x"0271",x"02BA",x"0004",x"0274",
    x"0298",x"0378",x"0020",x"0204",x"000C",x"02B8",x"0030",x"02B5",
    x"0274",x"0004",x"017C",x"039A",x"000C",x"000B",x"0012",x"022C",
    x"0010",x"02B4",x"02B1",x"0011",x"0065",x"0009",x"02B3",x"02B7",
    x"02B5",x"02B5",x"02B3",x"02B7",x"0275",x"0273",x"0271",x"008B",
    x"0274",x"02B4",x"0274",x"01C9",x"02A0",x"029D",x"037D",x"0020",
    x"0204",x"000B",x"0145",x"0204",x"0008",x"00D3",x"010B",x"029D",
    x"00AD",x"0204",x"0013",x"0220",x"0013",x"0009",x"014A",x"0204",
    x"0003",x"000B",x"0220",x"0017",x"02B4",x"00D4",x"0012",x"0113",
    x"0099",x"02B3",x"0119",x"0009",x"02B3",x"02B7",x"00A9",x"02B4",
    x"02B3",x"02B3",x"02B7",x"0275",x"02A0",x"0378",x"000D",x"0224",
    x"00DA",x"0081",x"03B9",x"00C0",x"0379",x"00C0",x"020C",x"0005",
    x"0014",x"0004",x"0128",x"02B2",x"02B7",x"0378",x"0041",x"022B",
    x"0014",x"0378",x"005B",x"0223",x"0018",x"0014",x"0004",x"0128",
    x"01B6",x"02B7",x"0275",x"02A0",x"0258",x"000B",x"02B8",x"0007",
    x"0040",x"0004",x"017C",x"039A",x"000C",x"0004",x"017C",x"039A",
    x"02A0",x"0014",x"0004",x"012C",x"01D2",x"0201",x"0004",x"0004",
    x"01E8",x"02F0",x"02B7",x"02B8",x"008B",x"0004",x"0128",x"01A8",
    x"02A0",x"0378",x"008C",x"0204",x"002F",x"0378",x"002E",x"0204",
    x"0013",x"0378",x"0085",x"020C",x"0006",x"0014",x"02B8",x"002D",
    x"0260",x"0200",x"0009",x"0378",x"002D",x"0204",x"0005",x"0004",
    x"012C",x"01D2",x"0201",x"0006",x"0014",x"0004",x"01E8",x"02F0",
    x"0200",x"000C",x"0378",x"0041",x"022B",x"0025",x"0378",x"005B",
    x"0223",x"0029",x"0014",x"0004",x"0128",x"01B6",x"02B8",x"008C",
    x"0004",x"0128",x"01A8",x"02B7",x"02B9",x"0041",x"0259",x"000B",
    x"0014",x"0220",x"000C",x"000A",x"037A",x"0007",x"020C",x"0095",
    x"0014",x"02B8",x"000D",x"0260",x"01C0",x"0260",x"02B3",x"02B4",
    x"00A2",x"02B7",x"0001",x"02F9",x"0004",x"0041",x"028B",x"00AF",
    x"0034",x"0034",x"0275",x"0001",x"02BA",x"0064",x"0001",x"0295",
    x"02FD",x"0200",x"02A8",x"0001",x"0378",x"0005",x"0023",x"0204",
    x"0017",x"0081",x"0001",x"03B9",x"0007",x"0036",x"0001",x"0379",
    x"0000",x"0022",x"0224",x"0011",x"0001",x"03B8",x"00F8",x"0009",
    x"0001",x"03F8",x"0000",x"0010",x"0015",x"0268",x"0220",x"001D",
    x"02B7",x"0046",x"004F",x"0052",x"0020",x"004E",x"0045",x"0058",
    x"0054",x"0052",x"0045",x"004D",x"0020",x"0044",x"0041",x"0054",
    x"0041",x"0044",x"0049",x"004D",x"0020",x"0049",x"0046",x"0020",
    x"0020",x"0050",x"0052",x"0049",x"004E",x"0045",x"004E",x"0044",
    x"0020",x"0047",x"004F",x"0054",x"004F",x"0047",x"0053",x"0055",
    x"0042",x"0043",x"004C",x"0052",x"0020",x"0049",x"004E",x"0050",
    x"0055",x"0052",x"0045",x"0054",x"0020",x"0043",x"0041",x"004C",
    x"004C",x"0053",x"0045",x"0054",x"0020",x"0050",x"0055",x"0054",
    x"0020",x"0047",x"0045",x"0054",x"0020",x"0052",x"0045",x"0041",
    x"0044",x"0049",x"0046",x"0020",x"0020",x"0000",x"003C",x"003D",
    x"003E",x"0028",x"002D",x"002B",x"002F",x"002A",x"00FF",x"0029",
    x"0275",x"0274",x"01D2",x"0273",x"01DB",x"02A0",x"0378",x"000D",
    x"0224",x"0093",x"0378",x"0022",x"020C",x"0002",x"03FB",x"0001",
    x"009B",x"022C",x"000D",x"0378",x"002C",x"020C",x"000A",x"0014",
    x"0004",x"0128",x"01A8",x"0014",x"02B8",x"000D",x"0260",x"0220",
    x"00B5",x"0001",x"02BD",x"0096",x"002B",x"0001",x"037D",x"00A0",
    x"002B",x"0224",x"0025",x"02A9",x"0141",x"022C",x"0009",x"0001",
    x"033D",x"0096",x"002B",x"03FD",x"0080",x"0014",x"0265",x"037D",
    x"0084",x"0224",x"0035",x"0220",x"00D1",x"0034",x"0275",x"0004",
    x"012C",x"03B7",x"0378",x"0022",x"020C",x"0022",x"0014",x"0004",
    x"0128",x"01A8",x"02A0",x"0378",x"0022",x"0204",x"0012",x"0378",
    x"000D",x"0204",x"0015",x"0258",x"000B",x"0001",x"02B8",x"0002",
    x"0006",x"0004",x"017C",x"039A",x"0012",x"0204",x"0016",x"0220",
    x"0016",x"0014",x"0004",x"0128",x"01A8",x"0004",x"012C",x"03B7",
    x"0378",x"002C",x"0204",x"000E",x"0378",x"000D",x"020C",x"0011",
    x"02A0",x"0080",x"0204",x"000C",x"0014",x"02B8",x"0001",x"0258",
    x"000B",x"02B7",x"0014",x"0004",x"0128",x"01A8",x"0220",x"000A",
    x"0014",x"0014",x"0220",x"000E",x"0275",x"02A0",x"0378",x"000D",
    x"0224",x"026B",x"0378",x"0041",x"022B",x"0008",x"0378",x"0044",
    x"0223",x"000C",x"0082",x"02B8",x"0124",x"0004",x"017C",x"039A",
    x"02A0",x"0378",x"000D",x"0224",x"027E",x"0378",x"0024",x"022C",
    x"0008",x"02B8",x"0124",x"0004",x"017C",x"039A",x"033A",x"0040",
    x"025A",x"000B",x"02B7",x"0275",x"0273",x"01DB",x"0004",x"0178",
    x"0252",x"009C",x"02B3",x"0224",x"0296",x"0011",x"00CF",x"0004",
    x"0128",x"02B2",x"02B7",x"0004",x"0128",x"01F2",x"02B7",x"0275",
    x"0280",x"015D",x"0081",x"03B9",x"0008",x"0204",x"006A",x"0081",
    x"03B9",x"0002",x"0204",x"0006",x"03B8",x"00F1",x"0240",x"015D",
    x"0200",x"012C",x"0081",x"03B9",x"0010",x"020C",x"0136",x"03B8",
    x"00F7",x"0240",x"015D",x"0283",x"0354",x"009C",x"02FC",x"002D",
    x"02A1",x"0379",x"00B0",x"020C",x"000A",x"02A1",x"0004",x"0120",
    x"03A3",x"009C",x"0004",x"0120",x"03AE",x"0200",x"0021",x"009C",
    x"0004",x"01E8",x"030C",x"0004",x"0174",x"01D4",x"0001",x"02B9",
    x"00FA",x"0047",x"028C",x"0001",x"02FC",x"00AF",x"0040",x"0014",
    x"00A2",x"0004",x"0178",x"008B",x"0281",x"035C",x"0004",x"01EC",
    x"0058",x"02FC",x"0002",x"02A0",x"0378",x"000D",x"020C",x"000F",
    x"0280",x"015D",x"03B8",x"0004",x"0204",x"00E1",x"02B8",x"0001",
    x"0001",x"02BD",x"0097",x"002D",x"0275",x"0200",x"017C",x"0001",
    x"033C",x"00AF",x"0040",x"0001",x"02B9",x"00FA",x"0047",x"024C",
    x"0280",x"015D",x"03B8",x"00E7",x"03F8",x"0018",x"0240",x"015D",
    x"02B7",x"0081",x"03B9",x"0004",x"020C",x"00B3",x"0081",x"03B9",
    x"0010",x"0204",x"0005",x"03B8",x"00FD",x"0240",x"015D",x"02B7",
    x"0001",x"02BD",x"00FC",x"0047",x"0001",x"02A9",x"008F",x"0284",
    x"0354",x"0004",x"012C",x"03B7",x"0378",x"000D",x"0204",x"00AE",
    x"0014",x"0001",x"02B9",x"009A",x"0026",x"02BA",x"0004",x"0004",
    x"0128",x"0264",x"0089",x"0204",x"0087",x"0011",x"0065",x"0009",
    x"00F9",x"02CF",x"006C",x"0058",x"0054",x"0074",x"007D",x"02B0",
    x"0065",x"0008",x"0004",x"012C",x"0274",x"03BA",x"0003",x"004E",
    x"004A",x"008D",x"00D7",x"0001",x"02BC",x"009A",x"0026",x"02BA",
    x"0004",x"0200",x"0016",x"0001",x"02BC",x"0049",x"002B",x"02BA",
    x"0004",x"0200",x"000E",x"0001",x"02BC",x"00EC",x"0026",x"02BA",
    x"0002",x"0200",x"0006",x"0001",x"02BC",x"00BB",x"0026",x"02BA",
    x"0004",x"0285",x"0354",x"00AB",x"02FB",x"000F",x"0091",x"02A0",
    x"0080",x"0204",x"000A",x"0268",x"0011",x"022C",x"0007",x"02B9",
    x"0020",x"0269",x"015D",x"022C",x"000E",x"02B9",x"000D",x"0269",
    x"0270",x"0272",x"0274",x"0004",x"012C",x"02DE",x"02B4",x"02B2",
    x"02B0",x"0080",x"022C",x"0022",x"0200",x"0041",x"02BA",x"0004",
    x"0200",x"000F",x"02BA",x"0002",x"0004",x"017C",x"00F0",x"0080",
    x"0204",x"0035",x"0004",x"012C",x"036C",x"0200",x"0030",x"02BA",
    x"0001",x"0004",x"017C",x"00F0",x"0200",x"0029",x"0004",x"012C",
    x"0274",x"0004",x"012C",x"01DE",x"0200",x"0021",x"0014",x"0004",
    x"012C",x"0274",x"0004",x"012C",x"028B",x"0200",x"0018",x"0004",
    x"0174",x"0212",x"0200",x"0013",x"0004",x"0124",x"0340",x"0200",
    x"000E",x"0081",x"03B9",x"0002",x"0204",x"0006",x"03B8",x"00F9",
    x"0240",x"015D",x"0200",x"000A",x"0004",x"012C",x"0224",x"0284",
    x"0354",x"02B8",x"006E",x"0004",x"0114",x"0338",x"0280",x"015D",
    x"0081",x"03B8",x"00EF",x"03B9",x"0004",x"020C",x"0004",x"03B8",
    x"00FD",x"03F8",x"0010",x"0240",x"015D",x"02B7",x"0275",x"01D2",
    x"02A0",x"0378",x"0020",x"0224",x"0004",x"0004",x"012C",x"01D2",
    x"0201",x"0016",x"0338",x"0030",x"0083",x"0090",x"02B9",x"000A",
    x"0004",x"011C",x"01DC",x"00DA",x"02B8",x"0322",x"0004",x"017C",
    x"039A",x"02A0",x"0001",x"037A",x"0080",x"000C",x"022B",x"001A",
    x"0014",x"02B7",x"0006",x"0378",x"0030",x"020B",x"0005",x"0378",
    x"003A",x"0203",x"0001",x"00AF",x"0007",x"00AF",x"0275",x"0004",
    x"0174",x"01F2",x"0092",x"020C",x"0005",x"009B",x"020C",x"0002",
    x"0013",x"0063",x"01E4",x"0280",x"015D",x"03B8",x"0002",x"020C",
    x"0032",x"0004",x"012C",x"020D",x"0004",x"012C",x"025A",x"0004",
    x"01E4",x"038F",x"02B4",x"0274",x"0004",x"0178",x"0320",x"03B9",
    x"0080",x"0204",x"0002",x"03F8",x"0007",x"0004",x"012C",x"02E9",
    x"0200",x"00CE",x"0034",x"0034",x"0034",x"0275",x"0004",x"01EC",
    x"039F",x"0048",x"0060",x"0204",x"000D",x"0150",x"022B",x"0009",
    x"0204",x"0003",x"0143",x"020B",x"0005",x"02B5",x"0272",x"0273",
    x"0274",x"00AF",x"02B5",x"02B7",x"0275",x"0280",x"0102",x"0378",
    x"0002",x"020D",x"0001",x"02B7",x"0001",x"02BD",x"00B5",x"0047",
    x"0001",x"02AC",x"00A4",x"0204",x"001E",x"0004",x"012C",x"025A",
    x"0004",x"0120",x"003B",x"0001",x"02BD",x"00B5",x"0047",x"0001",
    x"02AC",x"0080",x"0224",x"001E",x"020B",x"000D",x"0004",x"01EC",
    x"039F",x"022B",x"0004",x"0204",x"0006",x"01C0",x"0004",x"0120",
    x"0156",x"0220",x"002D",x"0280",x"015D",x"03B8",x"00FB",x"0240",
    x"015D",x"02B7",x"0275",x"0014",x"02A2",x"0285",x"0354",x"02FD",
    x"002A",x"00EA",x"033C",x"0003",x"02A0",x"0268",x"016A",x"022C",
    x"0004",x"01C0",x"0001",x"037D",x"00FA",x"0040",x"0204",x"0003",
    x"0268",x"0220",x"0008",x"02B7",x"0275",x"0004",x"012C",x"01AE",
    x"0272",x"0014",x"02A0",x"0378",x"000D",x"0204",x"0006",x"0378",
    x"002C",x"0204",x"0002",x"0220",x"000A",x"0004",x"012C",x"01AE",
    x"0093",x"02B2",x"02B7",x"0275",x"01E4",x"0004",x"012C",x"020D",
    x"0004",x"012C",x"0298",x"02B4",x"02B3",x"02B2",x"0220",x"000B",
    x"0275",x"00A5",x"033D",x"0002",x"02A8",x"03B8",x"0080",x"020C",
    x"0019",x"000D",x"02A8",x"0378",x"00A4",x"020C",x"0013",x"02A9",
    x"0339",x"00CB",x"0004",x"0128",x"031A",x"01C0",x"0248",x"0001",
    x"02BD",x"0009",x"0041",x"0001",x"02AA",x"004F",x"00DA",x"0004",
    x"012C",x"03BE",x"0014",x"02A0",x"033C",x"0003",x"0001",x"02BD",
    x"0007",x"0041",x"0275",x"0001",x"02A9",x"00A5",x"00C5",x"0169",
    x"0204",x"0004",x"02A8",x"0260",x"0220",x"0006",x"00A5",x"01C0",
    x"0268",x"0268",x"02B5",x"00A2",x"026A",x"0042",x"026A",x"02B7",
    x"02B4",x"02B3",x"02B2",x"0220",x"00F1",x"0034",x"0275",x"0001",
    x"02BD",x"00B3",x"0047",x"0001",x"02A8",x"0004",x"012C",x"02E9",
    x"02B7",x"0275",x"02BA",x"015E",x"0291",x"008B",x"03B9",x"0080",
    x"0204",x"000F",x"03BB",x"00BD",x"03FB",x"0040",x"0253",x"0291",
    x"03B9",x"0040",x"022C",x"0004",x"0291",x"03F9",x"0002",x"0251",
    x"02B7",x"0284",x"0354",x"02B5",x"0275",x"0270",x"0283",x"0163",
    x"02FB",x"0200",x"0004",x"01EC",x"0299",x"02B3",x"0282",x"0167",
    x"02FA",x"0200",x"0285",x"0163",x"0245",x"0164",x"02FD",x"0200",
    x"0155",x"020C",x"0013",x"0275",x"0274",x"0273",x"0272",x"0004",
    x"0178",x"03C7",x"0280",x"0164",x"0338",x"0014",x"0240",x"0164",
    x"02B2",x"02B3",x"02B4",x"02B5",x"033D",x"0014",x"02A1",x"0379",
    x"000D",x"0204",x"000B",x"0089",x"0204",x"0004",x"0339",x"0020",
    x"004D",x"0049",x"01D9",x"0269",x"0220",x"0025",x"0001",x"02B9",
    x"0005",x"0023",x"0269",x"033D",x"0200",x"0283",x"0164",x"011D",
    x"02FB",x"0014",x"033D",x"0015",x"020B",x"0002",x"02FB",x"0014",
    x"0243",x"0163",x"02FB",x"0200",x"0004",x"01EC",x"027E",x"02B7",
    x"0001",x"02BC",x"00B1",x"0047",x"0001",x"02B8",x"000A",x"0047",
    x"0260",x"0040",x"0260",x"0001",x"02B8",x"00E7",x"002C",x"02FC",
    x"0049",x"0260",x"0040",x"0260",x"0275",x"0004",x"012C",x"03ED",
    x"0001",x"02BD",x"00B1",x"0047",x"0275",x"0001",x"02A8",x"0270",
    x"0120",x"0004",x"0114",x"0338",x"0001",x"02BC",x"000D",x"0047",
    x"0274",x"02B8",x"00EF",x"0004",x"0114",x"0338",x"02B4",x"02B8",
    x"0040",x"0260",x"02FC",x"0003",x"0001",x"037C",x"005D",x"0047",
    x"022B",x"0008",x"0001",x"02BD",x"0007",x"0041",x"00A8",x"02F8",
    x"0004",x"0268",x"0040",x"0268",x"02B0",x"0268",x"0040",x"0268",
    x"02B5",x"0040",x"0268",x"0040",x"0268",x"0001",x"02B9",x"00B7",
    x"0047",x"02B8",x"0002",x"0248",x"0339",x"0003",x"02B8",x"0022",
    x"0248",x"02B7",x"0004",x"012C",x"036C",x"0220",x"021F",x"0275",
    x"02A0",x"0378",x"0020",x"0224",x"0004",x"02B7",x"0275",x"0001",
    x"02BD",x"0004",x"0041",x"02A9",x"004D",x"00CA",x"0001",x"037D",
    x"0007",x"0041",x"022C",x"0008",x"0001",x"02BD",x"0004",x"0041",
    x"0001",x"02BB",x"00FE",x"0040",x"02A9",x"004D",x"010A",x"000A",
    x"0090",x"0258",x"0040",x"000B",x"0258",x"000B",x"0012",x"0001",
    x"037D",x"0007",x"0041",x"022C",x"0010",x"0001",x"02BD",x"0009",
    x"0041",x"026A",x"0042",x"026A",x"02B7",x"0001",x"02BC",x"00CD",
    x"0047",x"0244",x"035C",x"0001",x"02BC",x"0085",x"0040",x"0244",
    x"0354",x"00AF",x"03FF",x"03FF",x"03FF",x"03FF",x"03FF",x"0021",
    x"0001",x"02B8",x"00C0",x"0007",x"0001",x"02BC",x"0040",x"0040",
    x"0004",x"0114",x"0338",x"0001",x"02BB",x"0051",x"002A",x"0001",
    x"02BA",x"00FF",x"002F",x"0253",x"0001",x"02BB",x"0001",x"00C0",
    x"0004",x"0120",x"001F",x"02A2",x"037A",x"01C1",x"020C",x"0003",
    x"0004",x"03C0",x"0043",x"0004",x"0320",x"0000",x"0001",x"02BB",
    x"0001",x"00E0",x"0004",x"0120",x"001F",x"0004",x"0110",x"00AB",
    x"000C",x"00A9",x"0041",x"03B9",x"00FD",x"0379",x"0001",x"0204",
    x"0006",x"0001",x"02B8",x"0023",x"0071",x"0240",x"02F0",x"0004",
    x"0310",x"003D",x"0002",x"0004",x"0114",x"00F1",x"0280",x"015E",
    x"0240",x"011E",x"0080",x"022C",x"000A",x"0001",x"02B8",x"0006",
    x"0019",x"0240",x"035D",x"0280",x"015F",x"0378",x"0002",x"020B",
    x"0061",x"020E",x"000C",x"0004",x"012C",x"0358",x"0001",x"02B8",
    x"0014",x"0050",x"0240",x"02F0",x"0004",x"0112",x"003D",x"0001",
    x"02B8",x"0098",x"0070",x"0240",x"035D",x"02B8",x"00E0",x"0240",
    x"015F",x"0004",x"0174",x"0052",x"0281",x"015F",x"03B9",x"0080",
    x"0204",x"0003",x"0004",x"0174",x"00DF",x"0200",x"004F",x"0275",
    x"0271",x"0281",x"035C",x"0004",x"01E0",x"02F5",x"004A",x"00D7",
    x"02B1",x"02B5",x"02B4",x"02B7",x"0378",x"002D",x"0204",x"0006",
    x"0378",x"0085",x"0204",x"0002",x"0006",x"00AF",x"0007",x"00AF",
    x"0052",x"0074",x"0065",x"0074",x"009A",x"0074",x"00AB",x"0074",
    x"0000",x"0000",x"0275",x"0281",x"035C",x"0004",x"01E0",x"02F5",
    x"01C0",x"0092",x"02B7",x"0034",x"0034",x"0034",x"0034",x"0034",
    x"0275",x"0281",x"00E0",x"02BD",x"000A",x"0015",x"022C",x"0002",
    x"007D",x"02B7",x"0004",x"012C",x"0358",x"0004",x"0174",x"01C7",
    x"02B8",x"0031",x"0240",x"015D",x"0001",x"02BD",x"0040",x"0040",
    x"0001",x"02A8",x"0080",x"0204",x"0001",x"0087",x"0004",x"0170",
    x"0251",x"0002",x"0280",x"0102",x"0010",x"0223",x"0005",x"0281",
    x"0103",x"0241",x"0102",x"0020",x"0004",x"0114",x"027D",x"0004",
    x"0114",x"00F1",x"0004",x"0110",x"01FA",x"0004",x"0114",x"03D5",
    x"0280",x"015E",x"0070",x"0209",x"0003",x"0004",x"0170",x"0134",
    x"0004",x"0118",x"02AD",x"0280",x"015D",x"03B8",x"0010",x"0204",
    x"0003",x"0004",x"01EC",x"00AC",x"0280",x"015D",x"0070",x"0209",
    x"0003",x"0004",x"012C",x"005F",x"0280",x"015F",x"03B8",x"0080",
    x"0204",x"0003",x"0004",x"0174",x"0117",x"0220",x"003D",x"00B5",
    x"0074",x"001B",x"0071",x"006F",x"0071",x"00D7",x"0074",x"0030",
    x"0071",x"002B",x"0071",x"0000",x"0000",x"0001",x"0001",x"0002",
    x"0003",x"0004",x"0005",x"0180",x"0190",x"01A0",x"01B0",x"01C0",
    x"01D0",x"01E0",x"01F0",x"0052",x"0045",x"0043",x"0053",x"0000",
    x"0002",x"0000",x"001B",x"0070",x"0275",x"0004",x"0170",x"015C",
    x"0280",x"015E",x"03B8",x"00DF",x"03F8",x"0020",x"0240",x"015E",
    x"02B9",x"011F",x"0282",x"00FF",x"03BA",x"00FF",x"0004",x"0114",
    x"012F",x"02B9",x"0120",x"0282",x"00FE",x"03BA",x"00FF",x"0004",
    x"0114",x"012F",x"0280",x"015E",x"03B8",x"00DF",x"0240",x"015E",
    x"0004",x"0170",x"015C",x"02B7",x"0275",x"02B8",x"0006",x"02BA",
    x"011F",x"0001",x"02BB",x"0042",x"0040",x"0294",x"029D",x"0255",
    x"025C",x"000A",x"000B",x"0010",x"022C",x"0008",x"02B7",x"0001",
    x"02BD",x"0042",x"0070",x"0275",x"02BA",x"0003",x"0242",x"00E0",
    x"0004",x"01EC",x"032B",x"02BB",x"00F0",x"0004",x"0174",x"01A0",
    x"0001",x"02B9",x"0049",x"0040",x"02B8",x"0023",x"0248",x"02B8",
    x"0080",x"0240",x"015E",x"0001",x"02B8",x"0085",x"0040",x"0001",
    x"02BC",x"004A",x"0040",x"0260",x"0040",x"0260",x"0004",x"0170",
    x"0213",x"0001",x"02B8",x"00C4",x"0071",x"0240",x"035D",x"02B7",
    x"0031",x"003A",x"0020",x"0042",x"0041",x"0053",x"0049",x"0043",
    x"0000",x"0029",x"0032",x"003A",x"0020",x"0043",x"0041",x"0052",
    x"0054",x"0052",x"0049",x"0044",x"0047",x"0045",x"0000",x"0051",
    x"0033",x"003A",x"0020",x"004D",x"0055",x"0053",x"0049",x"0043",
    x"0000",x"0079",x"0000",x"00FF",x"0000",x"0000",x"00CE",x"0071",
    x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0275",x"0081",
    x"0009",x"00F9",x"02CF",x"0024",x"002C",x"0032",x"0038",x"000C",
    x"000C",x"000C",x"0012",x"0012",x"0012",x"0025",x"004D",x"0082",
    x"0008",x"03B8",x"0003",x"0200",x"0005",x"0082",x"02F8",x"0021",
    x"03B8",x"0023",x"0001",x"02B9",x"0049",x"0040",x"0248",x"004E",
    x"004A",x"0001",x"03FA",x"0080",x"0022",x"0242",x"02AA",x"02B7",
    x"0004",x"0170",x"0213",x"01C0",x"0240",x"015F",x"02B7",x"0240",
    x"015F",x"02B9",x"0037",x"0200",x"000A",x"0240",x"015F",x"02B9",
    x"005F",x"0200",x"0004",x"0240",x"015F",x"02B9",x"0087",x"0004",
    x"0170",x"0224",x"02B7",x"0275",x"0001",x"02BB",x"0007",x"0022",
    x"0001",x"02B9",x"00A0",x"0071",x"0004",x"0170",x"0236",x"02B7",
    x"01C0",x"0240",x"015E",x"02B7",x"0001",x"02B8",x"0000",x"0022",
    x"0240",x"0237",x"0240",x"025F",x"0240",x"0287",x"02F9",x"0200",
    x"0001",x"02B8",x"0051",x"0022",x"0248",x"00AF",x"0275",x"0271",
    x"0004",x"0174",x"01C7",x"02B1",x"02BA",x"0200",x"008D",x"02A8",
    x"0080",x"022C",x"0003",x"02AC",x"037C",x"00FF",x"0204",x"0008",
    x"00D4",x"0004",x"0118",x"0067",x"00A9",x"0009",x"0220",x"0010",
    x"02B7",x"0275",x"0003",x"0001",x"02B8",x"0061",x"0000",x"0240",
    x"0100",x"0001",x"02B8",x"0072",x"0000",x"0240",x"0101",x"0002",
    x"02B7",x"0275",x"0004",x"0110",x"0126",x"0280",x"015D",x"03B8",
    x"0020",x"0204",x"0003",x"0004",x"0178",x"03E0",x"0280",x"015E",
    x"03B8",x"0008",x"0204",x"0003",x"0004",x"017C",x"0270",x"0280",
    x"015E",x"03B8",x"0040",x"0204",x"0003",x"0004",x"017C",x"03C0",
    x"0280",x"015F",x"03B8",x"0040",x"0204",x"0003",x"0004",x"0170",
    x"0293",x"0280",x"015F",x"03B8",x"0020",x"0204",x"0003",x"0004",
    x"0170",x"02B8",x"02B7",x"0275",x"0004",x"0174",x"005B",x"0001",
    x"02BB",x"004C",x"0040",x"009C",x"009D",x"02B8",x"0007",x"00C5",
    x"02A1",x"0269",x"0010",x"022C",x"0004",x"02B8",x"0040",x"0240",
    x"011E",x"02FB",x"0007",x"0018",x"02BC",x"00FE",x"0260",x"02A2",
    x"001A",x"0013",x"025A",x"0018",x"0060",x"022C",x"000B",x"02B7",
    x"0275",x"0004",x"0170",x"0318",x"0004",x"0170",x"02E0",x"02B7",
    x"0275",x"0001",x"02BB",x"004C",x"0040",x"00C3",x"029A",x"02FB",
    x"0007",x"029B",x"01D3",x"009B",x"02B7",x"0275",x"01C0",x"00A5",
    x"0001",x"02BC",x"005A",x"0040",x"0365",x"0204",x"0006",x"0008",
    x"0378",x"0006",x"022C",x"0007",x"02B7",x"0014",x"00A4",x"02B7",
    x"0275",x"01C0",x"0004",x"0170",x"02C0",x"0204",x"0028",x"01C9",
    x"007B",x"0209",x"001F",x"007A",x"0209",x"001D",x"0270",x"0272",
    x"0004",x"0170",x"035D",x"02BC",x"00FF",x"0004",x"0170",x"02CD",
    x"0204",x"001B",x"0262",x"0004",x"0170",x"034E",x"0280",x"015F",
    x"03B8",x"0080",x"0204",x"0002",x"0242",x"0169",x"02B2",x"02B0",
    x"0200",x"0001",x"0062",x"0009",x"009B",x"022C",x"0026",x"0008",
    x"0378",x"0007",x"022C",x"0031",x"02B7",x"02B2",x"02B0",x"02B7",
    x"0275",x"01C0",x"0004",x"0170",x"02C0",x"0204",x"0021",x"01C9",
    x"007B",x"0209",x"0018",x"007A",x"0201",x"0016",x"0270",x"0272",
    x"0004",x"0170",x"035D",x"0094",x"0004",x"0170",x"02CD",x"0204",
    x"0006",x"02BA",x"00FF",x"0262",x"0004",x"0170",x"0346",x"02B2",
    x"02B0",x"0200",x"0001",x"0062",x"0009",x"009B",x"022C",x"001F",
    x"0008",x"0378",x"0007",x"022C",x"002A",x"02B7",x"0275",x"0271",
    x"01C9",x"0004",x"0174",x"0163",x"02B1",x"02B7",x"0275",x"0271",
    x"0004",x"0170",x"0365",x"0004",x"0174",x"0153",x"02B9",x"000C",
    x"0004",x"0174",x"0163",x"02B1",x"02B7",x"0275",x"0082",x"004E",
    x"004A",x"00CA",x"02C2",x"0168",x"02B7",x"0275",x"0001",x"02BD",
    x"006F",x"0073",x"00D5",x"00D5",x"0001",x"02A9",x"02B7",x"005D",
    x"000D",x"009C",x"000C",x"00E7",x"000B",x"003C",x"000B",x"009B",
    x"000A",x"0002",x"000A",x"0073",x"0009",x"00EB",x"0008",x"006B",
    x"0008",x"00F2",x"0007",x"0080",x"0007",x"0014",x"0007",x"00AE",
    x"0006",x"004E",x"0006",x"00F4",x"0005",x"009E",x"0005",x"004D",
    x"0005",x"0001",x"0005",x"00B9",x"0004",x"0075",x"0004",x"0035",
    x"0004",x"00F9",x"0003",x"00C0",x"0003",x"008A",x"0003",x"0057",
    x"0003",x"0027",x"0003",x"00FA",x"0002",x"00CF",x"0002",x"00A7",
    x"0002",x"0081",x"0002",x"005D",x"0002",x"003B",x"0002",x"001B",
    x"0002",x"00FC",x"0001",x"00E0",x"0001",x"00C5",x"0001",x"00AC",
    x"0001",x"0094",x"0001",x"007D",x"0001",x"0068",x"0001",x"0053",
    x"0001",x"0040",x"0001",x"002E",x"0001",x"001D",x"0001",x"000D",
    x"0001",x"00FE",x"0000",x"00F0",x"0000",x"00E2",x"0000",x"00D6",
    x"0000",x"00CA",x"0000",x"00BE",x"0000",x"00B4",x"0000",x"00AA",
    x"0000",x"00A0",x"0000",x"0097",x"0000",x"008F",x"0000",x"0087",
    x"0000",x"007F",x"0000",x"0078",x"0000",x"0071",x"0000",x"006B",
    x"0000",x"0065",x"0000",x"005F",x"0000",x"005A",x"0000",x"0055",
    x"0000",x"0050",x"0000",x"004C",x"0000",x"0047",x"0000",x"0043",
    x"0000",x"0040",x"0000",x"003C",x"0000",x"0039",x"0000",x"0035",
    x"0000",x"0032",x"0000",x"0030",x"0000",x"002D",x"0000",x"002A",
    x"0000",x"0028",x"0000",x"0026",x"0000",x"0024",x"0000",x"0022",
    x"0000",x"0020",x"0000",x"001E",x"0000",x"001C",x"0000",x"001B",
    x"0000",x"0019",x"0000",x"0018",x"0000",x"0016",x"0000",x"0015",
    x"0000",x"0014",x"0000",x"0013",x"0000",x"0012",x"0000",x"0011",
    x"0000",x"0010",x"0000",x"000F",x"0000",x"000E",x"0000",x"0275",
    x"02B8",x"000E",x"0001",x"02BC",x"004C",x"0040",x"0004",x"0114",
    x"0338",x"02B8",x"0006",x"02B9",x"00FF",x"0001",x"02BC",x"005A",
    x"0040",x"0004",x"0114",x"0341",x"02BB",x"01F0",x"0004",x"0174",
    x"01A0",x"02BB",x"00F0",x"0004",x"0174",x"01A0",x"0004",x"0174",
    x"005B",x"02B7",x"0275",x"02B9",x"000C",x"0241",x"0168",x"0004",
    x"0174",x"002F",x"02B7",x"0275",x"02BB",x"00F8",x"0299",x"03B9",
    x"003F",x"03F9",x"0040",x"0259",x"02B7",x"0275",x"0378",x"0006",
    x"020E",x"002F",x"0281",x"0168",x"0048",x"00C7",x"0200",x"0029",
    x"0200",x"000A",x"0200",x"0025",x"0200",x"0009",x"0200",x"000A",
    x"0200",x"001F",x"0200",x"000A",x"0009",x"0200",x"000F",x"0011",
    x"0200",x"0006",x"02F9",x"000C",x"0200",x"0008",x"0339",x"000C",
    x"0089",x"0203",x"0009",x"01C9",x"0200",x"0006",x"0379",x"0030",
    x"0206",x"0002",x"02B9",x"0030",x"0241",x"0168",x"0004",x"0174",
    x"002F",x"02B7",x"0275",x"0080",x"020B",x"000C",x"0281",x"0168",
    x"0009",x"0379",x"0030",x"020D",x"0005",x"0241",x"0168",x"0004",
    x"0174",x"002F",x"02B7",x"0275",x"0080",x"022B",x"0004",x"0281",
    x"0168",x"0011",x"0223",x"000E",x"02B7",x"0001",x"0001",x"0001",
    x"0001",x"0001",x"0001",x"0001",x"0001",x"0001",x"0001",x"0001",
    x"0007",x"000F",x"000F",x"000E",x"0000",x"0001",x"0001",x"0001",
    x"0001",x"0001",x"0001",x"0011",x"0059",x"0071",x"00D9",x"0071",
    x"00D7",x"004F",x"000F",x"000E",x"0000",x"0000",x"0000",x"0000",
    x"0000",x"0000",x"00FF",x"0000",x"0000",x"0000",x"00FF",x"0275",
    x"02B8",x"00F0",x"02B9",x"0006",x"0041",x"02BC",x"0200",x"0004",
    x"0114",x"0341",x"02BC",x"023C",x"02B9",x"000E",x"0041",x"02B8",
    x"0064",x"0004",x"0114",x"0341",x"02BD",x"0264",x"02F9",x"0008",
    x"0261",x"0269",x"037C",x"02B4",x"022C",x"0005",x"0001",x"02B8",
    x"0041",x"0090",x"0001",x"02B9",x"00D4",x"0074",x"02BC",x"031D",
    x"02BA",x"00FF",x"0242",x"0169",x"0260",x"0261",x"0262",x"02FC",
    x"0005",x"037C",x"035D",x"022C",x"0008",x"0200",x"0037",x"0275",
    x"02B8",x"00FF",x"0283",x"0169",x"0143",x"0204",x"0033",x"0240",
    x"0169",x"0204",x"002F",x"0284",x"0324",x"0280",x"016A",x"02F8",
    x"0011",x"0240",x"016A",x"0078",x"02F8",x"000C",x"0040",x"0260",
    x"02B9",x"0069",x"0339",x"000E",x"033B",x"000C",x"022D",x"0005",
    x"02FB",x"0007",x"020B",x"0001",x"000B",x"02FB",x"0005",x"007B",
    x"01C0",x"0050",x"004B",x"0119",x"0041",x"0261",x"000C",x"0260",
    x"02FC",x"0004",x"037C",x"035F",x"020C",x"0002",x"02BC",x"031F",
    x"0244",x"0324",x"02B7",x"0275",x"0270",x"0273",x"0004",x"0174",
    x"0194",x"00C3",x"0259",x"0041",x"02FB",x"0004",x"0259",x"0041",
    x"02B3",x"02B0",x"02B7",x"0275",x"0270",x"0273",x"0004",x"0174",
    x"0194",x"02FB",x"000B",x"00C3",x"0259",x"02B3",x"02B0",x"02B7",
    x"0275",x"0270",x"0273",x"0274",x"0004",x"0174",x"0194",x"009C",
    x"02FC",x"0003",x"0262",x"0042",x"009C",x"02FC",x"0007",x"0262",
    x"0042",x"02FB",x"000A",x"0259",x"02B4",x"02B3",x"02B0",x"02B7",
    x"0275",x"0270",x"0273",x"0004",x"0174",x"0194",x"02FB",x"0009",
    x"0259",x"02B3",x"02B0",x"02B7",x"0378",x"0003",x"020B",x"0005",
    x"02BB",x"00F0",x"0338",x"0003",x"00AF",x"02BB",x"01F0",x"00AF",
    x"0275",x"0270",x"0273",x"0274",x"02B8",x"000E",x"009C",x"0004",
    x"0114",x"0338",x"02FB",x"0008",x"02B8",x"0038",x"0258",x"02B4",
    x"02B3",x"02B0",x"02B7",x"0275",x"0004",x"01EC",x"03B8",x"0284",
    x"0166",x"0280",x"0167",x"0120",x"02F8",x"0014",x"02FC",x"0200",
    x"02B9",x"0022",x"0041",x"0004",x"0114",x"0341",x"02B7",x"0275",
    x"0001",x"02B9",x"0000",x"0022",x"02BC",x"0200",x"02B8",x"00F0",
    x"0004",x"0114",x"0341",x"02B7",x"0275",x"0281",x"035C",x"02F9",
    x"0004",x"0288",x"03B8",x"0080",x"0204",x"0013",x"0339",x"0004",
    x"0288",x"0001",x"02BD",x"00D4",x"0047",x"00AB",x"0268",x"01C0",
    x"0268",x"0268",x"02B8",x"0001",x"0268",x"01C0",x"0004",x"01E0",
    x"0059",x"02B7",x"02B9",x"0011",x"0241",x"00E0",x"0001",x"02B9",
    x"0049",x"0040",x"0289",x"0241",x"00E2",x"01C0",x"0001",x"02B9",
    x"0048",x"0040",x"0248",x"00AF",x"00A3",x"0299",x"0379",x"00A0",
    x"020C",x"0007",x"0013",x"0299",x"0339",x"0008",x"00CB",x"01C9",
    x"0259",x"00AF",x"0275",x"01E4",x"02B9",x"00A0",x"0004",x"0174",
    x"02A1",x"0080",x"0204",x"000C",x"00A5",x"000D",x"02A9",x"02BB",
    x"00A1",x"01D2",x"00A0",x"0004",x"0174",x"02B0",x"0220",x"0013",
    x"01E4",x"02B9",x"00A1",x"0004",x"0174",x"02A1",x"0080",x"0204",
    x"000C",x"00A5",x"000D",x"02A9",x"02BB",x"00A0",x"0082",x"01C0",
    x"0004",x"0174",x"02B0",x"0220",x"0013",x"01E4",x"02B9",x"00A8",
    x"0004",x"0174",x"0322",x"02B9",x"00A9",x"0004",x"0174",x"0322",
    x"02B9",x"00B2",x"0004",x"0174",x"0322",x"01E4",x"0004",x"01EC",
    x"039F",x"0080",x"0204",x"000D",x"0223",x"0007",x"0082",x"004A",
    x"0062",x"01DB",x"0274",x"0004",x"012C",x"01DE",x"02B4",x"0220",
    x"0012",x"01E4",x"0004",x"01EC",x"039F",x"0080",x"0204",x"0022",
    x"022B",x"0007",x"00A3",x"0001",x"02BD",x"00B5",x"0047",x"026B",
    x"0043",x"026B",x"0004",x"0174",x"0204",x"0280",x"015D",x"03B8",
    x"00FB",x"03F8",x"0004",x"0240",x"015D",x"0001",x"02B9",x"00C2",
    x"0047",x"01C0",x"0248",x"01E4",x"0004",x"0174",x"028B",x"0004",
    x"0174",x"0292",x"02B7",x"0275",x"02B9",x"00A3",x"0004",x"0174",
    x"02A1",x"02B7",x"0275",x"0080",x"0204",x"0001",x"00A0",x"0001",
    x"02BD",x"00E9",x"0047",x"0268",x"0040",x"0268",x"01C0",x"0268",
    x"02B7",x"0275",x"0004",x"01EC",x"039F",x"022B",x"0004",x"0204",
    x"0005",x"00A5",x"02AA",x"014A",x"022C",x"000B",x"0080",x"02B7",
    x"0275",x"0274",x"0084",x"037B",x"00A0",x"020C",x"0002",x"01C0",
    x"0270",x"0004",x"01EC",x"039F",x"0080",x"022B",x"0005",x"0142",
    x"0204",x"0047",x"00A5",x"02A8",x"0158",x"0204",x"000E",x"037B",
    x"00A1",x"022C",x"0011",x"0378",x"00A0",x"022C",x"0015",x"02A8",
    x"0141",x"0204",x"0036",x"0220",x"001B",x"02A8",x"0141",x"022C",
    x"001F",x"037B",x"00A1",x"020C",x"0041",x"0274",x"0004",x"01EC",
    x"039F",x"0080",x"0204",x"0018",x"022B",x"0007",x"00A5",x"02A8",
    x"02AA",x"0378",x"00A0",x"020C",x"0003",x"0151",x"0204",x"000C",
    x"0378",x"00A1",x"022C",x"0015",x"0151",x"022C",x"0018",x"0004",
    x"0174",x"0314",x"0220",x"001D",x"02B4",x"00A0",x"02B4",x"00A5",
    x"0015",x"02A9",x"0339",x"0005",x"00CD",x"0268",x"0040",x"0268",
    x"02B7",x"037B",x"00A0",x"020C",x"0004",x"02B4",x"00A4",x"022C",
    x"0013",x"02B4",x"0200",x"0001",x"0275",x"00A5",x"033D",x"0002",
    x"02A8",x"03F8",x"0080",x"0015",x"0268",x"02B7",x"02B5",x"0274",
    x"0220",x"0068",x"0275",x"01E4",x"0271",x"02B1",x"0271",x"0004",
    x"0174",x"02A1",x"0204",x"001D",x"0274",x"00A5",x"0015",x"02A9",
    x"00CD",x"033D",x"0005",x"0001",x"02AA",x"01E4",x"0004",x"01EC",
    x"039F",x"0204",x"0006",x"0142",x"022C",x"0007",x"02B4",x"0220",
    x"001B",x"02B4",x"0004",x"0174",x"0314",x"02B5",x"02B5",x"0220",
    x"010B",x"02B5",x"02B7",x"0275",x"00A2",x"033A",x"0006",x"0001",
    x"037A",x"00AF",x"0040",x"0204",x"0005",x"0290",x"0378",x"0080",
    x"0224",x"000C",x"02FA",x"0005",x"0290",x"0378",x"0082",x"0204",
    x"0008",x"0378",x"000D",x"0204",x"0004",x"0378",x"0001",x"022C",
    x"001B",x"0095",x"000D",x"01C9",x"008A",x"0090",x"02AB",x"037B",
    x"0080",x"020C",x"000D",x"02AB",x"009B",x"0204",x"0005",x"0091",
    x"00AA",x"0012",x"0012",x"0008",x"02FD",x"0004",x"0200",x"0027",
    x"03BB",x"00C0",x"037B",x"00C0",x"020C",x"000D",x"0091",x"00AA",
    x"0012",x"0008",x"02AB",x"037B",x"0080",x"020C",x"0012",x"02FD",
    x"0005",x"0200",x"000E",x"0015",x"02AB",x"037B",x"0041",x"020B",
    x"0008",x"037B",x"005B",x"0203",x"0004",x"0091",x"00AA",x"0012",
    x"0008",x"02AB",x"037B",x"002D",x"0204",x"0001",x"0015",x"016C",
    x"022C",x"003B",x"0092",x"020C",x"0001",x"008A",x"0378",x"0002",
    x"020B",x"0020",x"02B8",x"0002",x"0093",x"0004",x"0178",x"00D8",
    x"015C",x"0204",x"0005",x"0010",x"0020",x"0094",x"0010",x"02B7",
    x"008B",x"0004",x"0178",x"00D8",x"015A",x"0204",x"0001",x"0010",
    x"0080",x"0224",x"000C",x"0378",x"0002",x"022C",x"0011",x"008C",
    x"0220",x"0013",x"0378",x"0001",x"022C",x"000D",x"0093",x"0004",
    x"0178",x"00D8",x"015C",x"0224",x"0014",x"0220",x"0022",x"0275",
    x"00A5",x"01C0",x"02A9",x"0379",x"000D",x"0204",x"0011",x"0379",
    x"0080",x"020C",x"0004",x"02FD",x"0005",x"0220",x"000C",x"03B9",
    x"00E0",x"0379",x"0080",x"022C",x"0012",x"0008",x"0015",x"00AC",
    x"02B7",x"0275",x"02A0",x"0378",x"0080",x"020C",x"0007",x"01C0",
    x"0260",x"00A2",x"02FC",x"0004",x"0200",x"004B",x"0081",x"03B8",
    x"00C0",x"0378",x"00C0",x"020C",x"003C",x"0014",x"01C0",x"0260",
    x"02A0",x"0378",x"0080",x"020C",x"002B",x"01C0",x"0260",x"00A2",
    x"02FC",x"0004",x"0274",x"02B8",x"0001",x"0270",x"03B9",x"003F",
    x"02BB",x"0016",x"02B8",x"0008",x"0004",x"01EC",x"03E0",x"0159",
    x"020B",x"0009",x"0119",x"0285",x"02F0",x"02FD",x"000A",x"0001",
    x"02AC",x"0200",x"0004",x"0001",x"02BC",x"006E",x"0026",x"0049",
    x"00CC",x"0001",x"02A3",x"02B0",x"009F",x"02B4",x"0200",x"0011",
    x"0014",x"00A2",x"0004",x"0178",x"008B",x"01C0",x"0260",x"0220",
    x"002E",x"00A2",x"0012",x"0093",x"0004",x"0178",x"008B",x"01C0",
    x"0258",x"02A0",x"0378",x"002D",x"020C",x"001D",x"0095",x"000D",
    x"00A9",x"02F9",x"0003",x"02A8",x"0080",x"020C",x"0005",x"0169",
    x"022C",x"0006",x"0200",x"000F",x"0091",x"0001",x"02BA",x"00DB",
    x"0047",x"0004",x"01EC",x"0058",x"033A",x"0004",x"0291",x"03F9",
    x"0080",x"0251",x"000C",x"0014",x"02A0",x"0080",x"0224",x"0003",
    x"0378",x"000D",x"0204",x"000D",x"0378",x"0080",x"020C",x"0009",
    x"02A0",x"0080",x"020C",x"0004",x"02FC",x"0004",x"0220",x"0013",
    x"0014",x"0014",x"02B7",x"0275",x"0292",x"033A",x"0041",x"004E",
    x"0001",x"02FA",x"000D",x"0047",x"02B7",x"0275",x"03BA",x"001F",
    x"033A",x"0005",x"000A",x"00FA",x"02D7",x"0004",x"0009",x"000C",
    x"000F",x"02B8",x"0001",x"0004",x"03E0",x"005A",x"01C0",x"0220",
    x"0005",x"0004",x"03E0",x"0268",x"0004",x"03E0",x"00BC",x"0275",
    x"0001",x"02BC",x"00B2",x"0040",x"02A0",x"03B8",x"00C0",x"0378",
    x"00C0",x"0204",x"000A",x"0014",x"0004",x"0174",x"03F9",x"0281",
    x"035C",x"0004",x"01EC",x"0058",x"02B7",x"00A2",x"0014",x"0291",
    x"0379",x"0080",x"020C",x"0004",x"02FA",x"0002",x"0200",x"0003",
    x"0004",x"0178",x"008B",x"02A1",x"01C0",x"0270",x"0220",x"00B9",
    x"0275",x"009D",x"02AB",x"037B",x"0080",x"020C",x"0004",x"02FD",
    x"0005",x"0200",x"0013",x"03BB",x"00C0",x"037B",x"00C0",x"020C",
    x"0007",x"02AB",x"037B",x"0080",x"020C",x"0002",x"02FD",x"0005",
    x"02AB",x"037B",x"002D",x"0204",x"0001",x"0015",x"00AB",x"02B7",
    x"0275",x"0001",x"02BA",x"00EE",x"0047",x"02A0",x"0378",x"000D",
    x"0204",x"00AF",x"0378",x"002D",x"0204",x"001D",x"0081",x"03B9",
    x"00F0",x"0379",x"0080",x"0204",x"0064",x"0081",x"03B9",x"00C0",
    x"0379",x"00C0",x"0204",x"0043",x"0378",x"002E",x"0204",x"0005",
    x"0004",x"012C",x"01D2",x"0201",x"0014",x"0014",x"0004",x"01E8",
    x"02F0",x"0220",x"0025",x"02A0",x"0014",x"0378",x"002E",x"0224",
    x"000B",x"0004",x"012C",x"01D2",x"0229",x"0010",x"000C",x"0220",
    x"002A",x"0378",x"0041",x"022B",x"0037",x"0378",x"005B",x"0223",
    x"003B",x"033C",x"0002",x"02A0",x"0270",x"0378",x"002D",x"020C",
    x"0005",x"02B8",x"0032",x"0004",x"017C",x"039A",x"02A0",x"0258",
    x"000B",x"02B8",x"0024",x"0004",x"017C",x"039A",x"02B0",x"0378",
    x"002D",x"022C",x"0055",x"0258",x"000B",x"0220",x"0059",x"033C",
    x"0002",x"02A0",x"0378",x"002D",x"020C",x"000E",x"02B8",x"0032",
    x"0004",x"017C",x"039A",x"0004",x"0128",x"02B2",x"02B8",x"002D",
    x"0258",x"000B",x"0220",x"006E",x"0004",x"0128",x"02B2",x"0220",
    x"0073",x"0001",x"02B8",x"0026",x"0005",x"0004",x"017C",x"039A",
    x"0014",x"02A0",x"0378",x"0084",x"020C",x"0004",x"0258",x"000B",
    x"0200",x"0025",x"0378",x"008A",x"020C",x"0011",x"0291",x"0379",
    x"0084",x"0204",x"0005",x"0259",x"000B",x"0012",x"0220",x"0009",
    x"02B9",x"008A",x"0259",x"000B",x"0012",x"0220",x"0099",x"0001",
    x"037A",x"00EE",x"0047",x"0204",x"000A",x"0291",x"0270",x"0008",
    x"0009",x"0060",x"0061",x"0148",x"02B0",x"0206",x"0004",x"000A",
    x"0250",x"0220",x"00AD",x"0291",x"0259",x"000B",x"0012",x"0220",
    x"0019",x"0001",x"037A",x"00EE",x"0047",x"0204",x"0006",x"0290",
    x"0258",x"000B",x"0012",x"0220",x"000B",x"02B7",x"0275",x"0273",
    x"0004",x"0178",x"020D",x"0094",x"01DB",x"0004",x"0178",x"0252",
    x"0204",x"0038",x"0004",x"0178",x"02CE",x"0204",x"0038",x"020B",
    x"000F",x"02BB",x"0001",x"0004",x"0178",x"0252",x"020E",x"0008",
    x"020B",x"000B",x"0014",x"02B8",x"0020",x"0260",x"0220",x"001C",
    x"0004",x"0178",x"02CE",x"0220",x"0017",x"0004",x"0178",x"0252",
    x"0204",x"0004",x"0223",x"000B",x"022B",x"0008",x"0014",x"02B8",
    x"0020",x"0260",x"00A5",x"02A8",x"0378",x"000D",x"0224",x"0034",
    x"0378",x"008A",x"022C",x"0008",x"0015",x"02B8",x"0020",x"0268",
    x"0220",x"003E",x"01C0",x"0010",x"02B3",x"0094",x"02B7",x"0004",
    x"0178",x"02F6",x"01C0",x"0220",x"0008",x"0275",x"00A2",x"0094",
    x"01C9",x"02A0",x"0378",x"000D",x"0204",x"0016",x"0378",x"0084",
    x"0204",x"0006",x"0378",x"008A",x"0204",x"0005",x"0220",x"000E",
    x"0009",x"0220",x"0011",x"0011",x"0223",x"0014",x"0014",x"02B8",
    x"0020",x"0260",x"0220",x"001C",x"0089",x"0204",x"000F",x"0094",
    x"02A0",x"0378",x"0084",x"022C",x"0004",x"02B8",x"0020",x"0014",
    x"0260",x"0011",x"022C",x"000B",x"0220",x"002E",x"02B7",x"0204",
    x"000C",x"0004",x"012C",x"01D2",x"0209",x"0007",x"0378",x"0045",
    x"020C",x"0005",x"01ED",x"000D",x"02B7",x"01ED",x"02B7",x"01ED",
    x"0015",x"02B7",x"0275",x"0272",x"0274",x"00A2",x"02A0",x"0378",
    x"000D",x"0204",x"006F",x"0378",x"0084",x"020C",x"0008",x"009B",
    x"0224",x"000C",x"02B5",x"02B2",x"01C9",x"0011",x"02B7",x"0378",
    x"0085",x"020C",x"0005",x"0014",x"02B8",x"002D",x"0260",x"02A0",
    x"0081",x"03B9",x"00C0",x"0379",x"00C0",x"020C",x"002B",x"000C",
    x"02A0",x"0004",x"012C",x"01D2",x"0209",x"002D",x"0014",x"02A0",
    x"0378",x"008B",x"022C",x"0004",x"02A0",x"0014",x"0378",x"0085",
    x"020C",x"0003",x"02B8",x"002D",x"0260",x"02A0",x"0378",x"008C",
    x"022C",x"0004",x"0093",x"02B5",x"02B2",x"0298",x"02B9",x"0001",
    x"03B8",x"00C0",x"0378",x"00C0",x"0204",x"0002",x"02F9",x"0004",
    x"0089",x"02B7",x"0378",x"002E",x"0204",x"0005",x"0004",x"012C",
    x"01D2",x"0201",x"0008",x"0004",x"01EC",x"003F",x"0223",x"0004",
    x"0014",x"0220",x"0020",x"0378",x"0041",x"020B",x"0006",x"0378",
    x"005B",x"0203",x"0002",x"0220",x"002A",x"033C",x"0002",x"02A0",
    x"0378",x"002D",x"020C",x"0001",x"0014",x"02B8",x"0020",x"0260",
    x"0220",x"0074",x"02B4",x"02B2",x"0200",x"0025",x"0275",x"00A5",
    x"02A8",x"0378",x"000D",x"0204",x"001E",x"0378",x"0085",x"020B",
    x"0008",x"0378",x"008A",x"0203",x"0004",x"00AC",x"01C9",x"0009",
    x"02B7",x"0378",x"008A",x"020C",x"0004",x"00AC",x"01C9",x"0011",
    x"02B7",x"0378",x"0084",x"0224",x"001C",x"02B8",x"0020",x"0015",
    x"0268",x"0220",x"0022",x"01C9",x"0089",x"02B7",x"0275",x"0094",
    x"02A0",x"0378",x"000D",x"0204",x"002E",x"0378",x"0084",x"022C",
    x"0008",x"00A5",x"02A8",x"0378",x"0020",x"0224",x"0004",x"0378",
    x"008A",x"0204",x"000D",x"0378",x"0085",x"022B",x"0016",x"0378",
    x"008A",x"0223",x"001A",x"02A8",x"0378",x"008A",x"022C",x"0004",
    x"0014",x"0015",x"02B8",x"0020",x"0260",x"0268",x"0220",x"0028",
    x"033C",x"0002",x"02A1",x"02B8",x"0022",x"0040",x"00AF",x"02B5",
    x"02B5",x"02B4",x"00A2",x"02B7",x"0275",x"0274",x"01D2",x"02A0",
    x"0378",x"000D",x"0224",x"000A",x"0378",x"0022",x"020C",x"0002",
    x"03FA",x"0001",x"0092",x"022C",x"000D",x"0014",x"02BA",x"002C",
    x"01C0",x"0004",x"01EC",x"03E0",x"0272",x"0200",x"0036",x"008D",
    x"02FD",x"0010",x"0001",x"02A9",x"02BA",x"0002",x"0004",x"0128",
    x"0264",x"02B2",x"00D1",x"0151",x"020C",x"000F",x"0001",x"02B9",
    x"00EC",x"0026",x"02BA",x"0002",x"0004",x"0128",x"0264",x"0089",
    x"020C",x"0003",x"000C",x"0220",x"0036",x"0274",x"0271",x"02A0",
    x"0004",x"012C",x"01D2",x"0201",x"0018",x"0274",x"02B2",x"02B1",
    x"02B4",x"0011",x"0061",x"03F9",x"00C0",x"033C",x"0002",x"0261",
    x"0261",x"0094",x"0220",x"004D",x"0034",x"0004",x"0120",x"002F",
    x"022E",x"003A",x"02B5",x"0220",x"002E",x"0014",x"02A0",x"0378",
    x"000D",x"0224",x"0063",x"0378",x"0084",x"022C",x"0008",x"0014",
    x"02B8",x"008B",x"0260",x"02A0",x"0378",x"000D",x"0224",x"0070",
    x"0378",x"0084",x"020C",x"0004",x"0014",x"02B8",x"0020",x"0260",
    x"0378",x"008A",x"022C",x"0010",x"0014",x"02B8",x"008C",x"0260",
    x"0274",x"0220",x"003C",x"0275",x"0001",x"02B8",x"0060",x"0040",
    x"0285",x"0160",x"00AA",x"03BD",x"000F",x"0066",x"0066",x"0155",
    x"020C",x"0002",x"01C9",x"02B7",x"00C5",x"02A9",x"0105",x"03BD",
    x"000F",x"004E",x"004E",x"00EA",x"0242",x"0160",x"02B7",x"0275",
    x"0284",x"0166",x"02FC",x"0200",x"00A5",x"02FD",x"0014",x"0282",
    x"0167",x"02FA",x"0200",x"02AB",x"0263",x"016A",x"022D",x"0004",
    x"02BB",x"0022",x"0043",x"0263",x"0162",x"022D",x"0003",x"02B7",
    x"0275",x"0004",x"0170",x"0293",x"0001",x"02BD",x"004C",x"0040",
    x"00AB",x"029A",x"0091",x"03BA",x"0080",x"01D1",x"0259",x"02FB",
    x"0007",x"0299",x"03B9",x"007F",x"0259",x"02FB",x"0005",x"0299",
    x"03B9",x"00BF",x"0259",x"033B",x"0007",x"0299",x"008C",x"03B9",
    x"0040",x"01CC",x"025C",x"01CA",x"000B",x"0299",x"01D1",x"0259",
    x"02B8",x"00FF",x"00B9",x"02F9",x"0011",x"033B",x"0006",x"009C",
    x"02A2",x"02FD",x"0007",x"0092",x"020C",x"0067",x"02F9",x"0008",
    x"02A2",x"016C",x"0225",x"0008",x"02B7",x"0008",x"002E",x"003B",
    x"0070",x"001B",x"0030",x"000D",x"0000",x"002C",x"006D",x"006B",
    x"0069",x"0039",x"0038",x"006F",x"006C",x"006E",x"0062",x"0068",
    x"0079",x"0037",x"0036",x"0075",x"006A",x"0076",x"0063",x"0066",
    x"0072",x"0035",x"0034",x"0074",x"0067",x"0078",x"007A",x"0073",
    x"0077",x"0033",x"0032",x"0065",x"0064",x"0020",x"000A",x"000B",
    x"0071",x"0031",x"000C",x"0000",x"0061",x"0025",x"003E",x"003A",
    x"0050",x"001B",x"0029",x"000D",x"0000",x"003C",x"004D",x"004B",
    x"0049",x"0028",x"002A",x"004F",x"004C",x"004E",x"0042",x"0048",
    x"0059",x"002F",x"002D",x"0055",x"004A",x"0056",x"0043",x"0046",
    x"0052",x"002B",x"0024",x"0054",x"0047",x"0058",x"005A",x"0053",
    x"0057",x"0023",x"0022",x"0045",x"0044",x"0020",x"003F",x"005E",
    x"0051",x"003D",x"0027",x"0000",x"0041",x"02FC",x"0006",x"02A3",
    x"0183",x"0204",x"0001",x"02B7",x"0006",x"0009",x"007A",x"0229",
    x"0003",x"0015",x"02AA",x"03BA",x"0080",x"0204",x"0002",x"02F9",
    x"0030",x"00CB",x"0299",x"0089",x"0204",x"0059",x"0015",x"02AA",
    x"03BA",x"0040",x"0204",x"000A",x"0379",x"0060",x"0205",x"0006",
    x"0379",x"007F",x"020E",x"0002",x"0339",x"0060",x"02BD",x"0019",
    x"0245",x"011E",x"0280",x"015E",x"0082",x"03B8",x"0010",x"0204",
    x"0005",x"01C2",x"0242",x"015E",x"0241",x"0161",x"0379",x"001B",
    x"020C",x"001D",x"0280",x"015D",x"03B8",x"00FD",x"02F8",x"0002",
    x"0240",x"015D",x"02BB",x"015E",x"0298",x"0081",x"03B9",x"0040",
    x"0204",x"0004",x"02B9",x"000D",x"0241",x"00E1",x"03B8",x"00B5",
    x"03F8",x"0002",x"0258",x"0004",x"0174",x"01F2",x"02B7",x"0280",
    x"0160",x"0082",x"03B8",x"000F",x"0066",x"0066",x"0093",x"000A",
    x"03BA",x"000F",x"0150",x"0204",x"000A",x"0001",x"02FB",x"0060",
    x"0040",x"0259",x"004E",x"004E",x"00D0",x"0240",x"0160",x"02B7",
    x"0275",x"0280",x"015E",x"03B8",x"003F",x"0240",x"015E",x"0280",
    x"015F",x"03B8",x"00E0",x"01D0",x"0240",x"015F",x"03B8",x"0004",
    x"020C",x"0006",x"0001",x"02BD",x"0080",x"0040",x"0200",x"0004",
    x"0001",x"02BD",x"00FA",x"0040",x"02B8",x"0020",x"02B9",x"0004",
    x"0268",x"0011",x"022C",x"0003",x"02A0",x"0378",x"0020",x"0224",
    x"0004",x"033D",x"0004",x"02B9",x"0004",x"0378",x"000D",x"0204",
    x"0005",x"0268",x"02A0",x"0011",x"022C",x"0008",x"0001",x"02BC",
    x"0085",x"0040",x"02B8",x"0041",x"0260",x"0001",x"037C",x"0089",
    x"0040",x"022C",x"0006",x"02B8",x"000D",x"0260",x"0004",x"012C",
    x"02DE",x"02B8",x"001D",x"0240",x"00E2",x"01C0",x"0004",x"017C",
    x"01DA",x"0004",x"017C",x"020D",x"01C0",x"0240",x"00E2",x"02B8",
    x"0005",x"0004",x"017C",x"01DA",x"0004",x"017C",x"020D",x"02B8",
    x"0005",x"0281",x"015F",x"02F8",x"0005",x"0079",x"0229",x"0004",
    x"0004",x"017C",x"01DA",x"0001",x"02B8",x"00FA",x"0040",x"0001",
    x"02BD",x"0007",x"0041",x"0001",x"02A9",x"02F9",x"0002",x"0282",
    x"015F",x"007E",x"0201",x"0007",x"0202",x"000A",x"0004",x"017C",
    x"0228",x"0200",x"000F",x"0004",x"017C",x"021C",x"0200",x"000A",
    x"0001",x"02BD",x"00B1",x"0047",x"0001",x"02A9",x"0009",x"0004",
    x"017C",x"0221",x"0280",x"015E",x"007C",x"0202",x"004B",x"007C",
    x"0222",x"0007",x"0280",x"015F",x"03B8",x"0004",x"0204",x"0001",
    x"02B7",x"0001",x"02B9",x"007B",x"0040",x"0001",x"02BB",x"0000",
    x"0022",x"0284",x"0163",x"02FC",x"01FA",x"0004",x"0118",x"0067",
    x"0280",x"015F",x"03B8",x"0010",x"0204",x"0011",x"00A3",x"02B9",
    x"0004",x"0013",x"0298",x"0001",x"03B8",x"00FF",x"0009",x"0001",
    x"03F8",x"0000",x"0010",x"0258",x"0011",x"022C",x"000D",x"0001",
    x"02BC",x"007B",x"0040",x"0001",x"02BD",x"0080",x"0040",x"02A8",
    x"0378",x"0020",x"0204",x"0008",x"0015",x"02A8",x"0360",x"022C",
    x"006D",x"0080",x"022C",x"0006",x"0280",x"015F",x"03B8",x"0010",
    x"0204",x"0007",x"0285",x"0163",x"033D",x"0014",x"0004",x"0328",
    x"0328",x"02B7",x"0275",x"0001",x"02BB",x"0006",x"0022",x"0001",
    x"02B9",x"00F4",x"007D",x"00C1",x"0284",x"0163",x"037C",x"0013",
    x"020E",x"0004",x"02FC",x"0014",x"0244",x"0163",x"02FC",x"01EC",
    x"0004",x"0118",x"0067",x"02B7",x"0053",x"0045",x"0054",x"0020",
    x"0000",x"0047",x"004F",x"0020",x"0020",x"0000",x"0056",x"0045",
    x"0052",x"0046",x"0000",x"004C",x"004F",x"0041",x"0044",x"0000",
    x"0053",x"0041",x"0056",x"0045",x"0000",x"0275",x"02BA",x"01FE",
    x"02BB",x"01FF",x"0004",x"0114",x"00B7",x"0290",x"0040",x"03D8",
    x"0018",x"0224",x"0005",x"02B7",x"0275",x"02BA",x"0107",x"0200",
    x"0003",x"0275",x"02BA",x"0207",x"02BB",x"001D",x"0200",x"0009",
    x"0275",x"0010",x"0011",x"0001",x"02BA",x"0000",x"0004",x"02BB",
    x"0039",x"0243",x"00E2",x"02BB",x"001D",x"0243",x"00E0",x"0001",
    x"02BC",x"0071",x"0040",x"0262",x"0042",x"0283",x"015F",x"03BB",
    x"00E0",x"01D3",x"0243",x"015F",x"0260",x"0040",x"0260",x"0261",
    x"0041",x"0261",x"0040",x"0041",x"0108",x"0260",x"0040",x"0260",
    x"02FC",x"0002",x"01C0",x"0260",x"02FC",x"0004",x"0260",x"02FC",
    x"0004",x"0260",x"0281",x"015E",x"03B9",x"00F5",x"03F9",x"0008",
    x"0241",x"015E",x"02B7",x"001E",x"0024",x"002E",x"0046",x"0047",
    x"0056",x"006C",x"007A",x"007D",x"0093",x"009F",x"00A8",x"00B5",
    x"0275",x"0001",x"02BB",x"0071",x"0040",x"0298",x"009A",x"0012",
    x"01C9",x"0001",x"02BC",x"0063",x"007E",x"00A5",x"00C4",x"02E5",
    x"00AF",x"02B9",x"0050",x"0251",x"0008",x"0258",x"02B7",x"0291",
    x"0011",x"0251",x"022C",x"0005",x"02B9",x"0049",x"0251",x"0220",
    x"000C",x"0281",x"00E0",x"007D",x"022A",x"000F",x"0291",x"0011",
    x"0251",x"0204",x"000A",x"03B9",x"0007",x"0204",x"0001",x"02B7",
    x"02B9",x"00AA",x"0241",x"00E1",x"02B7",x"0241",x"00E1",x"0220",
    x"0024",x"0011",x"0285",x"00E0",x"03BD",x"0002",x"0224",x"0029",
    x"009C",x"00CC",x"02FC",x"0006",x"02A1",x"0241",x"00E1",x"0220",
    x"0034",x"0281",x"00E0",x"007D",x"022A",x"0037",x"009C",x"000C",
    x"0004",x"017C",x"0362",x"028D",x"0245",x"00E1",x"0001",x"0361",
    x"022C",x"0043",x"02B9",x"0028",x"0251",x"0220",x"004A",x"0291",
    x"0011",x"0251",x"022C",x"004D",x"0241",x"00E2",x"0281",x"015E",
    x"03B9",x"00F7",x"0241",x"015E",x"02B7",x"0008",x"0200",x"0011",
    x"0004",x"0170",x"00B0",x"0229",x"005E",x"0281",x"00E1",x"0379",
    x"00AA",x"020C",x"0006",x"0291",x"0011",x"0251",x"0224",x"006B",
    x"02B7",x"02B9",x"0005",x"0251",x"0220",x"0070",x"0004",x"0170",
    x"00B0",x"0229",x"0074",x"0281",x"00E1",x"0379",x"00AA",x"022C",
    x"007C",x"02B7",x"0004",x"0170",x"00B0",x"0229",x"0080",x"02BC",
    x"0005",x"0200",x"0007",x"0004",x"0170",x"00B0",x"0229",x"0089",
    x"02BC",x"0006",x"00DC",x"0281",x"00E1",x"0261",x"0220",x"0093",
    x"0004",x"0170",x"00B0",x"0229",x"0096",x"03B9",x"0038",x"0204",
    x"0003",x"0004",x"017C",x"036E",x"009C",x"000C",x"0004",x"017C",
    x"0362",x"008A",x"0012",x"0281",x"00E1",x"02FB",x"0009",x"029D",
    x"037D",x"0004",x"020D",x"000E",x"000D",x"025D",x"0001",x"02FD",
    x"007A",x"0040",x"0269",x"0285",x"015F",x"03BD",x"0002",x"0204",
    x"0010",x"0251",x"0285",x"015F",x"03BD",x"0001",x"0204",x"0008",
    x"0351",x"0204",x"0006",x"0004",x"017C",x"036E",x"0200",x"0001",
    x"0251",x"033B",x"0009",x"0001",x"0362",x"0204",x"0006",x"0004",
    x"017C",x"0362",x"0224",x"0087",x"02B7",x"0004",x"017C",x"036E",
    x"0220",x"008D",x"0275",x"0001",x"02A1",x"0009",x"0014",x"0014",
    x"0261",x"0041",x"0261",x"0041",x"0089",x"02B7",x"0275",x"0281",
    x"015F",x"03B9",x"00EF",x"03F9",x"0010",x"0241",x"015F",x"02B7",
    x"0275",x"02A0",x"0378",x"0001",x"0204",x"001B",x"02B8",x"0022",
    x"0258",x"000B",x"0014",x"02A0",x"0378",x"0001",x"0204",x"0004",
    x"0258",x"000B",x"0220",x"0008",x"02B8",x"0022",x"0258",x"000B",
    x"02A0",x"0080",x"0204",x"0004",x"02B8",x"002C",x"0258",x"000B",
    x"0014",x"02B7",x"0275",x"0040",x"0281",x"0164",x"02F9",x"0200",
    x"00A5",x"0001",x"033D",x"0086",x"0040",x"00E9",x"028D",x"0001",
    x"03BD",x"00FF",x"0009",x"01C5",x"024D",x"0040",x"02B7",x"02A0",
    x"0080",x"020C",x"0003",x"0004",x"03E8",x"02DF",x"0275",x"02F8",
    x"0040",x"0258",x"000B",x"02B8",x"0024",x"0258",x"000B",x"02B7",
    x"0001",x"02B9",x"0049",x"0040",x"0289",x"03B9",x"0020",x"0204",
    x"002F",x"0280",x"00E0",x"03B8",x"000A",x"0378",x"0002",x"020C",
    x"0026",x"0001",x"02BC",x"004A",x"0040",x"0001",x"02A2",x"0001",
    x"02B9",x"0048",x"0040",x"028B",x"00DA",x"0292",x"0092",x"020C",
    x"0002",x"03FA",x"0020",x"0242",x"00E1",x"000B",x"024B",x"037A",
    x"000D",x"020C",x"000C",x"0281",x"015E",x"03B9",x"00BF",x"0241",
    x"015E",x"0001",x"02B9",x"0048",x"0040",x"01C0",x"0248",x"00AF",
    x"0281",x"00E0",x"03B9",x"0002",x"022C",x"002C",x"00AF",x"0170",
    x"0275",x"0285",x"0354",x"02FD",x"002A",x"0001",x"02A9",x"0049",
    x"0061",x"01E4",x"0004",x"01EC",x"039F",x"0048",x"0060",x"0204",
    x"0008",x"0141",x"022C",x"0009",x"0271",x"0004",x"012C",x"0298",
    x"02B1",x"01E4",x"0004",x"01EC",x"039F",x"0048",x"0060",x"0204",
    x"0003",x"0148",x"022B",x"0009",x"033C",x"0004",x"0001",x"02BD",
    x"0007",x"0041",x"0275",x"0001",x"02AA",x"0093",x"0001",x"02B9",
    x"00B1",x"0040",x"0289",x"00CB",x"0001",x"02A8",x"02B5",x"0143",
    x"020B",x"0003",x"0004",x"0328",x"0323",x"026B",x"0043",x"026B",
    x"0043",x"009D",x"01C0",x"0268",x"0268",x"0290",x"0258",x"0012",
    x"0013",x"0154",x"022C",x"0006",x"000C",x"0001",x"02BD",x"00AF",
    x"0040",x"00AB",x"00CB",x"02A8",x"0260",x"016B",x"022C",x"0004",
    x"02B7",x"0275",x"0274",x"0270",x"0004",x"01E0",x"0123",x"02B0",
    x"0080",x"0204",x"0004",x"0288",x"03F8",x"0080",x"0248",x"01C0",
    x"0001",x"02BB",x"00D4",x"0047",x"009C",x"033C",x"0007",x"0004",
    x"01E0",x"0147",x"0080",x"0204",x"000C",x"00A1",x"0080",x"020B",
    x"0002",x"02F9",x"0007",x"01C0",x"0004",x"01E0",x"015E",x"0220",
    x"0019",x"0004",x"01E0",x"0183",x"009B",x"0204",x"000A",x"0288",
    x"03B8",x"0080",x"020C",x"0002",x"0339",x"0007",x"0004",x"01E0",
    x"0194",x"0004",x"01E0",x"01C0",x"0004",x"01E0",x"0183",x"0339",
    x"0007",x"009B",x"020C",x"0008",x"0080",x"0204",x"0017",x"0004",
    x"01E0",x"015E",x"0200",x"0012",x"0080",x"020C",x"000B",x"0004",
    x"01E0",x"0194",x"028A",x"03BA",x"007F",x"03FA",x"0080",x"024A",
    x"0200",x"0004",x"028A",x"03BA",x"007F",x"024A",x"0004",x"01E0",
    x"021A",x"02B4",x"02B7",x"0275",x"0274",x"0284",x"035C",x"000C",
    x"00A5",x"02FD",x"0006",x"00A9",x"0298",x"0268",x"02A0",x"0268",
    x"014C",x"022C",x"0004",x"01C0",x"033C",x"0006",x"0260",x"014C",
    x"022C",x"0003",x"000B",x"009D",x"02FD",x"0003",x"0281",x"015D",
    x"03B9",x"0080",x"0204",x"0002",x"02FD",x"0003",x"02B9",x"0080",
    x"00AC",x"0098",x"0271",x"0004",x"01E0",x"01FD",x"00A5",x"0083",
    x"02B1",x"0298",x"0188",x"0204",x"0009",x"0275",x"0273",x"0271",
    x"0004",x"01E0",x"01C0",x"02B1",x"02B3",x"02B5",x"0061",x"0089",
    x"022C",x"0019",x"000B",x"015D",x"022C",x"001F",x"01C0",x"0270",
    x"0004",x"01E0",x"021A",x"0092",x"0204",x"01EC",x"0004",x"01E0",
    x"01DD",x"0093",x"02F9",x"0007",x"0004",x"01E0",x"01DD",x"02B0",
    x"0270",x"0080",x"0203",x"0001",x"0022",x"00DA",x"0339",x"0007",
    x"0004",x"01E0",x"01EB",x"0004",x"01E0",x"0183",x"0339",x"0007",
    x"028A",x"0200",x"01C7",x"0275",x"0272",x"0001",x"02BA",x"00D4",
    x"0047",x"0272",x"0153",x"0204",x"0017",x"0001",x"02B9",x"00FE",
    x"0025",x"0004",x"01EC",x"005C",x"033A",x"0007",x"02B8",x"0004",
    x"0281",x"015D",x"03B9",x"0080",x"0204",x"0002",x"02F8",x"0003",
    x"0099",x"0004",x"01EC",x"005E",x"02B1",x"02B2",x"02B7",x"0275",
    x"0099",x"0004",x"01E0",x"01DD",x"0090",x"00A1",x"0004",x"01E0",
    x"01DD",x"0142",x"0204",x"0005",x"020B",x"0005",x"02B8",x"0001",
    x"02B7",x"01C0",x"02B7",x"01C0",x"0010",x"02B7",x"0275",x"0004",
    x"01E0",x"01DD",x"000A",x"0004",x"01E0",x"01EB",x"0082",x"004E",
    x"004E",x"0090",x"008A",x"02F9",x"0007",x"000A",x"0151",x"0204",
    x"000F",x"0293",x"009D",x"0067",x"0067",x"01C3",x"0253",x"03BD",
    x"000F",x"00AB",x"004F",x"004F",x"0098",x"000A",x"0220",x"0011",
    x"0339",x"0007",x"02B7",x"0275",x"0281",x"035C",x"028A",x"02F9",
    x"0007",x"028D",x"03BA",x"0080",x"03BD",x"0080",x"01DB",x"0155",
    x"0204",x"0001",x"000B",x"02B7",x"0275",x"0004",x"01E0",x"02F5",
    x"0092",x"020C",x"0005",x"028A",x"03BA",x"007F",x"024A",x"02B7",
    x"008C",x"0009",x"02FC",x"0007",x"028B",x"001B",x"03BB",x"00FF",
    x"024B",x"0009",x"014C",x"022C",x"0008",x"0011",x"033C",x"0007",
    x"02BB",x"0001",x"028A",x"00DA",x"0093",x"03BA",x"00FF",x"024A",
    x"0043",x"03BB",x"00FF",x"0011",x"014C",x"022C",x"000C",x"02B7",
    x"01C0",x"0001",x"02B9",x"00D3",x"0047",x"008A",x"02FA",x"0007",
    x"028B",x"0294",x"00E3",x"00C3",x"009C",x"03BC",x"00FF",x"024C",
    x"0043",x"03BB",x"00FF",x"0098",x"0011",x"0012",x"0001",x"037A",
    x"00D4",x"0047",x"022C",x"0013",x"00AF",x"0275",x"028A",x"03BA",
    x"007F",x"0095",x"03BD",x"0040",x"020C",x"0002",x"0022",x"02B7",
    x"03FA",x"0040",x"02B7",x"0275",x"0092",x"0203",x"0003",x"0022",
    x"0200",x"0002",x"03FA",x"0040",x"028D",x"03BD",x"0080",x"0204",
    x"0002",x"03FA",x"0080",x"024A",x"02B7",x"0275",x"0001",x"02B9",
    x"00D5",x"0047",x"01ED",x"028A",x"0062",x"01EA",x"0095",x"028A",
    x"024D",x"03BA",x"0001",x"0204",x"0004",x"02BD",x"0080",x"0200",
    x"0001",x"01ED",x"0009",x"0001",x"0379",x"00DB",x"0047",x"022C",
    x"0015",x"02B7",x"0275",x"0281",x"035C",x"0004",x"01E0",x"02F5",
    x"0092",x"020C",x"0004",x"02B8",x"0040",x"0248",x"02B7",x"0009",
    x"028A",x"03BA",x"00F0",x"020C",x"0022",x"0011",x"0004",x"01E0",
    x"01DD",x"0012",x"0004",x"01E0",x"01EB",x"02F9",x"0006",x"01E4",
    x"028A",x"0095",x"03BA",x"000F",x"004E",x"004E",x"01E2",x"024A",
    x"00AA",x"03BA",x"00F0",x"0066",x"0066",x"0094",x"0011",x"0001",
    x"0379",x"00CD",x"0047",x"022C",x"0014",x"0220",x"0027",x"0011",
    x"02B7",x"0275",x"009D",x"00C5",x"000C",x"000B",x"015D",x"0224",
    x"00FF",x"0298",x"02A1",x"0148",x"0224",x"0008",x"0148",x"020B",
    x"0003",x"02B8",x"0001",x"02B7",x"01C0",x"0010",x"02B7",x"0275",
    x"0274",x"0004",x"01E0",x"0123",x"008C",x"02B8",x"0007",x"00C4",
    x"0004",x"0114",x"0338",x"0004",x"01E0",x"02F5",x"0092",x"020C",
    x"0007",x"0004",x"011C",x"031D",x"02B4",x"0004",x"03EC",x"004A",
    x"0004",x"0170",x"007F",x"0034",x"00A3",x"02B8",x"0007",x"0103",
    x"0004",x"01E0",x"0251",x"0080",x"020B",x"0006",x"0281",x"035C",
    x"01C0",x"0004",x"01E0",x"015E",x"02B8",x"0080",x"0001",x"02BB",
    x"00DB",x"0047",x"0004",x"01E0",x"01FD",x"009A",x"008B",x"033B",
    x"000E",x"009C",x"0270",x"02B8",x"0007",x"00C4",x"0004",x"01E0",
    x"0251",x"0083",x"02B0",x"009B",x"020B",x"001B",x"0291",x"01C1",
    x"0251",x"0272",x"0270",x"0001",x"02B9",x"00D4",x"0047",x"0004",
    x"01E0",x"02F5",x"0092",x"0204",x"000A",x"0004",x"01E0",x"0194",
    x"0004",x"01E0",x"01C0",x"0091",x"0004",x"01E0",x"0194",x"02B0",
    x"02B2",x"0093",x"0060",x"022C",x"0032",x"000B",x"02B8",x"0080",
    x"0001",x"037B",x"00E1",x"0047",x"022C",x"003B",x"0284",x"035C",
    x"000C",x"00A5",x"02FD",x"000D",x"00A1",x"02F9",x"0006",x"02A8",
    x"0260",x"0161",x"022C",x"0004",x"0339",x"0007",x"01C0",x"0010",
    x"0220",x"01EA",x"03BA",x"007F",x"009B",x"0204",x"0002",x"03FA",
    x"0080",x"024A",x"02B4",x"02B4",x"02B7",x"0275",x"008D",x"02F9",
    x"0007",x"000D",x"02AA",x"0092",x"020C",x"0005",x"0169",x"022C",
    x"0006",x"0200",x"0002",x"02BA",x"0001",x"0339",x"0007",x"02B7",
    x"0275",x"0004",x"01EC",x"0049",x"0091",x"0282",x"035C",x"0004",
    x"01EC",x"0058",x"02B8",x"0001",x"0004",x"01E0",x"0059",x"01C0",
    x"0281",x"035C",x"0004",x"01E0",x"02F5",x"0092",x"0204",x"000A",
    x"0284",x"035C",x"02A1",x"03B9",x"0080",x"0008",x"0089",x"0204",
    x"0001",x"0020",x"02B7",x"0004",x"01E0",x"03BD",x"0004",x"01E4",
    x"0000",x"0004",x"01E4",x"0019",x"02B5",x"02B5",x"02B5",x"0200",
    x"0152",x"0004",x"01E0",x"03BD",x"0004",x"01E0",x"03E6",x"0220",
    x"000F",x"0004",x"01E0",x"03BD",x"0004",x"01E4",x"0000",x"0004",
    x"01E4",x"0029",x"0004",x"01E4",x"002E",x"0220",x"001A",x"0004",
    x"01E0",x"03BD",x"0004",x"01E0",x"03E6",x"0220",x"000F",x"0001",
    x"02B9",x"0051",x"0047",x"008B",x"033B",x"0028",x"0288",x"02BC",
    x"011F",x"03B8",x"0080",x"0204",x"0001",x"000C",x"02A0",x"0081",
    x"0082",x"03B8",x"000F",x"03B9",x"0040",x"0204",x"0002",x"02F8",
    x"0064",x"03BA",x"0080",x"020C",x"0002",x"0008",x"0020",x"0004",
    x"01E4",x"01FB",x"033B",x"001C",x"000C",x"02A0",x"0081",x"03B8",
    x"0003",x"0200",x"014B",x"02BB",x"0030",x"02BA",x"0007",x"0004",
    x"01E4",x"037D",x"0270",x"02BB",x"0034",x"0004",x"01E4",x"037D",
    x"0004",x"0114",x"0372",x"03BB",x"007F",x"02B0",x"0272",x"0273",
    x"0004",x"0114",x"0372",x"03BB",x"007F",x"02B1",x"0119",x"0203",
    x"0001",x"0021",x"02B0",x"0110",x"0203",x"0001",x"0020",x"00C8",
    x"0001",x"02BB",x"0019",x"0047",x"0200",x"0120",x"01C0",x"0270",
    x"0004",x"01E0",x"03C6",x"02B5",x"02B5",x"02B5",x"02B0",x"0008",
    x"0378",x"0006",x"022C",x"000C",x"02B7",x"0275",x"02BB",x"0008",
    x"02BA",x"0005",x"0004",x"01E4",x"037D",x"02B5",x"0275",x"0270",
    x"0004",x"0174",x"0194",x"02FB",x"0008",x"0084",x"0004",x"0114",
    x"0345",x"0082",x"0048",x"004C",x"01D0",x"029D",x"0018",x"0185",
    x"0018",x"01C5",x"025D",x"00DC",x"02FC",x"0003",x"01C0",x"0260",
    x"02B0",x"02B4",x"0273",x"0272",x"0270",x"00A7",x"0275",x"02BA",
    x"001F",x"02BB",x"003C",x"0004",x"01E4",x"037D",x"02B4",x"0081",
    x"02B0",x"0270",x"0004",x"0174",x"0188",x"02B0",x"02B2",x"02B3",
    x"029D",x"0091",x"0049",x"004D",x"01CD",x"025D",x"0220",x"001D",
    x"0275",x"0001",x"02BA",x"00FF",x"000F",x"02BB",x"003C",x"0004",
    x"01E4",x"037D",x"02B4",x"0081",x"02B0",x"0270",x"0004",x"0174",
    x"0153",x"02B0",x"02B2",x"02B3",x"0299",x"01D1",x"0259",x"0220",
    x"0036",x"0275",x"02BA",x"000F",x"02BB",x"0054",x"0004",x"01E4",
    x"037D",x"02B4",x"0081",x"02B0",x"0270",x"0004",x"0174",x"0163",
    x"00A7",x"0275",x"02B8",x"0030",x"0220",x"000C",x"0275",x"0001",
    x"02BB",x"0039",x"0047",x"0004",x"01E4",x"01A2",x"0270",x"02BB",
    x"0010",x"02BA",x"000F",x"0004",x"01E4",x"037D",x"0081",x"02B2",
    x"02B4",x"02B0",x"0270",x"0004",x"0174",x"0170",x"00A7",x"0001",
    x"02BB",x"0045",x"0047",x"02BC",x"0007",x"0004",x"01E4",x"01DC",
    x"0080",x"0203",x"0006",x"0020",x"0004",x"0114",x"02D5",x"0200",
    x"0032",x"0004",x"0114",x"02CF",x"0200",x"002D",x"0001",x"02BC",
    x"005D",x"0047",x"02B9",x"0001",x"0004",x"01EC",x"03CA",x"0004",
    x"01EC",x"0372",x"0274",x"02BB",x"0038",x"02BA",x"0007",x"0004",
    x"01E4",x"037D",x"0004",x"0114",x"036C",x"008A",x"02B1",x"0001",
    x"02BD",x"0000",x"0050",x"02AB",x"0043",x"03BB",x"00FC",x"020C",
    x"0020",x"02FD",x"0013",x"0245",x"02F0",x"0004",x"0114",x"02B2",
    x"0004",x"012C",x"03ED",x"02B8",x"0001",x"02B7",x"0001",x"02BD",
    x"0007",x"0041",x"0001",x"02A9",x"0001",x"02AA",x"0001",x"02BC",
    x"00B1",x"0047",x"0001",x"02A3",x"033A",x"0008",x"0151",x"020B",
    x"0005",x"0004",x"011C",x"031B",x"0220",x"001A",x"033B",x"0008",
    x"0273",x"033C",x"0002",x"0263",x"0043",x"0263",x"0004",x"012C",
    x"03BE",x"02BB",x"0030",x"02BA",x"000F",x"0004",x"01E4",x"037D",
    x"0008",x"0081",x"02B4",x"000C",x"0220",x"0059",x"02BB",x"0034",
    x"02BA",x"005F",x"0004",x"01E4",x"037D",x"0082",x"0004",x"0170",
    x"0365",x"0088",x"0001",x"02BB",x"0049",x"0047",x"0004",x"01EC",
    x"0340",x"0220",x"0047",x"0061",x"0339",x"0012",x"0004",x"0120",
    x"03A3",x"0270",x"0271",x"0093",x"02BA",x"0014",x"02B9",x"0001",
    x"0004",x"01E4",x"0191",x"02B1",x"00C1",x"0011",x"02B0",x"0080",
    x"020C",x"000B",x"0271",x"02BA",x"003F",x"0004",x"01E4",x"0387",
    x"02B1",x"02F8",x"0020",x"0248",x"02B7",x"0288",x"0080",x"0204",
    x"013B",x"0338",x"0020",x"0200",x"0137",x"0004",x"01E4",x"02B3",
    x"01C9",x"0200",x"0005",x"0004",x"01E4",x"02B3",x"02B9",x"0001",
    x"02FA",x"0004",x"0080",x"020C",x"001D",x"0271",x"0272",x"0283",
    x"035C",x"02BC",x"007F",x"0004",x"01E4",x"01DC",x"02B2",x"02B3",
    x"0270",x"0290",x"0004",x"0114",x"0357",x"02B5",x"009B",x"020C",
    x"0003",x"00A8",x"0200",x"0001",x"00A9",x"0004",x"0114",x"034F",
    x"0250",x"02B7",x"0290",x"008B",x"0004",x"0114",x"0357",x"009B",
    x"0204",x"003C",x"0088",x"0200",x"0039",x"0270",x"0093",x"0004",
    x"01E4",x"01A2",x"0378",x"0004",x"020C",x"001D",x"0001",x"02BD",
    x"00B3",x"0047",x"02B0",x"0080",x"0204",x"0006",x"0001",x"02A8",
    x"03B8",x"0007",x"0200",x"00E8",x"0275",x"02BA",x"0007",x"0004",
    x"01E4",x"0387",x"0001",x"03F8",x"0000",x"0022",x"02B5",x"0268",
    x"0040",x"0268",x"02B7",x"02B1",x"0089",x"0204",x"001C",x"0001",
    x"02BA",x"00B7",x"0047",x"0293",x"0063",x"0067",x"03BB",x"0003",
    x"0143",x"020C",x"000C",x"0290",x"03B8",x"0007",x"0001",x"02BB",
    x"00DB",x"0047",x"0004",x"01E4",x"01FB",x"0200",x"00C4",x"01C0",
    x"0010",x"0220",x"000C",x"0270",x"02BA",x"0007",x"0004",x"01E4",
    x"0387",x"02B1",x"0379",x"0004",x"020B",x"0002",x"02B9",x"0003",
    x"004D",x"0049",x"01C8",x"0001",x"02BA",x"00B7",x"0047",x"0250",
    x"02B7",x"0275",x"0271",x"0272",x"0004",x"01E4",x"01A2",x"02B2",
    x"02B1",x"0148",x"0203",x"0001",x"0088",x"0142",x"0203",x"0001",
    x"0090",x"02B7",x"0275",x"0099",x"0001",x"02BA",x"00DB",x"0047",
    x"0004",x"01EC",x"0058",x"0001",x"02BB",x"00DB",x"0047",x"0004",
    x"01E4",x"01B3",x"02B7",x"0275",x"0299",x"03B9",x"0080",x"020C",
    x"001E",x"0099",x"0004",x"01E0",x"01DD",x"0092",x"020B",x"0017",
    x"037A",x"0005",x"0203",x"0015",x"037A",x"0004",x"0204",x"0009",
    x"01C0",x"0004",x"01E0",x"015E",x"0004",x"01E0",x"01DD",x"0220",
    x"000C",x"008D",x"000D",x"0001",x"02A8",x"0040",x"02B7",x"01C0",
    x"02B7",x"01C0",x"0010",x"02B7",x"0275",x"0099",x"0001",x"02BA",
    x"00DB",x"0047",x"0093",x"0004",x"01EC",x"0058",x"0298",x"0081",
    x"03B9",x"0080",x"03B8",x"007F",x"0258",x"0271",x"0004",x"01E4",
    x"01B3",x"0144",x"0203",x"0001",x"00A0",x"02B5",x"00AD",x"0204",
    x"0001",x"0020",x"02B7",x"0275",x"01ED",x"0080",x"0203",x"0002",
    x"000D",x"0020",x"0275",x"0004",x"01EC",x"0340",x"02B5",x"00AD",
    x"0204",x"0004",x"0298",x"03F8",x"0080",x"0258",x"02B7",x"0004",
    x"01E4",x"02B3",x"02B9",x"00A7",x"0200",x"0006",x"0004",x"01E4",
    x"02B3",x"02B9",x"0068",x"000A",x"02FA",x"0002",x"0080",x"020C",
    x"0009",x"0272",x"008A",x"0004",x"01E4",x"0387",x"0040",x"02B2",
    x"0250",x"02B7",x"0290",x"0040",x"02BB",x"00FF",x"0379",x"00A7",
    x"0204",x"0001",x"0063",x"0198",x"0001",x"02BB",x"00DB",x"0047",
    x"0004",x"01EC",x"0340",x"009A",x"0004",x"0378",x"003D",x"0004",
    x"01E4",x"02B3",x"0272",x"0080",x"020C",x"0017",x"02BA",x"000F",
    x"0004",x"01E4",x"0387",x"02B2",x"0291",x"0001",x"03B9",x"00E8",
    x"00FF",x"0083",x"03B8",x"0007",x"03BB",x"0008",x"0204",x"0002",
    x"03F8",x"0010",x"01C1",x"0251",x"02B7",x"02B2",x"0294",x"00A5",
    x"03BD",x"0010",x"03BC",x"0007",x"00AD",x"0204",x"0002",x"03FC",
    x"0008",x"00A0",x"0220",x"0037",x"0080",x"0224",x"00CD",x"02B8",
    x"0064",x"0004",x"0114",x"029E",x"0220",x"0041",x"02BB",x"0010",
    x"0043",x"0273",x"0200",x"0000",x"0004",x"01E4",x"02B3",x"0272",
    x"0080",x"020C",x"0013",x"0283",x"035C",x"02B2",x"02B1",x"0019",
    x"0294",x"0298",x"03B8",x"0080",x"0204",x"0003",x"018C",x"0254",
    x"02B7",x"018C",x"0019",x"01CC",x"0254",x"02B7",x"02B2",x"02B1",
    x"0294",x"018C",x"00A4",x"0204",x"0002",x"02BC",x"0002",x"00A0",
    x"0010",x"0220",x"0134",x"02BB",x"0020",x"0220",x"002E",x"02BB",
    x"0001",x"0220",x"0032",x"02BB",x"0004",x"0220",x"0036",x"02BB",
    x"0002",x"0220",x"003A",x"0275",x"0270",x"0093",x"01C9",x"02BA",
    x"0007",x"0004",x"01E4",x"0191",x"0004",x"0114",x"036C",x"008A",
    x"02B0",x"02B7",x"0270",x"0061",x"0271",x"0001",x"02F9",x"00F9",
    x"0040",x"0288",x"0080",x"0204",x"0022",x"0270",x"0093",x"0004",
    x"01E4",x"01A2",x"02B1",x"0141",x"020B",x"0019",x"0080",x"0204",
    x"0016",x"02B2",x"004A",x"0095",x"0001",x"02FD",x"00E8",x"0040",
    x"0001",x"02AA",x"0010",x"004C",x"00C2",x"02B0",x"0080",x"022C",
    x"00AC",x"0281",x"035C",x"0004",x"01EC",x"0058",x"02B7",x"02B5",
    x"02B5",x"00AD",x"0224",x"0005",x"0001",x"02BA",x"00FE",x"0025",
    x"0220",x"00BD",x"0080",x"0224",x"000E",x"0093",x"0001",x"02BC",
    x"00FF",x"007F",x"0004",x"01E4",x"01DC",x"0220",x"0198",x"0270",
    x"0093",x"01C9",x"02BA",x"00EF",x"0004",x"01E4",x"0191",x"0081",
    x"02F9",x"0200",x"02B0",x"0080",x"020C",x"001B",x"0271",x"02BA",
    x"000F",x"0004",x"01E4",x"0387",x"0081",x"0082",x"03B8",x"0003",
    x"03B9",x"0004",x"03BA",x"0008",x"004A",x"004D",x"0049",x"0048",
    x"01C8",x"01D0",x"0040",x"02B1",x"0248",x"0004",x"01EC",x"03B8",
    x"02B7",x"028A",x"0042",x"0090",x"0091",x"03B8",x"0020",x"03B9",
    x"0010",x"03BA",x"0006",x"0062",x"0061",x"0064",x"0060",x"01C8",
    x"01D0",x"0220",x"010E",x"0004",x"01E4",x"02B3",x"02FA",x"0005",
    x"0080",x"020C",x"000F",x"0272",x"02BA",x"000F",x"0004",x"01E4",
    x"0387",x"02B2",x"0291",x"0001",x"03B9",x"00F0",x"00FF",x"01C1",
    x"0251",x"02B7",x"0290",x"03B8",x"000F",x"0220",x"012A",x"0004",
    x"01E4",x"02B3",x"02FA",x"0005",x"0080",x"020C",x"000F",x"0272",
    x"02BA",x"003F",x"0004",x"01E4",x"0387",x"02B2",x"0291",x"03B9",
    x"000F",x"004C",x"004C",x"01C1",x"0251",x"02B7",x"0290",x"0064",
    x"0064",x"03B8",x"003F",x"0220",x"0148",x"0275",x"0001",x"02FB",
    x"000D",x"0047",x"01C9",x"0004",x"01E4",x"0191",x"02B7",x"0275",
    x"0283",x"035C",x"01C9",x"0004",x"01E4",x"0191",x"02B7",x"0275",
    x"0284",x"0354",x"0274",x"02B8",x"0029",x"0004",x"0114",x"0338",
    x"02B3",x"009C",x"02FC",x"002A",x"0004",x"01E8",x"016B",x"000C",
    x"02B8",x"0012",x"0004",x"01EC",x"03E0",x"009D",x"02A1",x"0089",
    x"0204",x"0335",x"0088",x"03B8",x"00E0",x"0378",x"00A0",x"020C",
    x"010D",x"03B9",x"001F",x"004D",x"008A",x"0001",x"02FA",x"0049",
    x"002B",x"02BB",x"0004",x"0290",x"0378",x"0020",x"0204",x"0005",
    x"0268",x"000A",x"0013",x"022C",x"0009",x"02B8",x"0020",x"0268",
    x"00AB",x"0065",x"0009",x"00F9",x"02CF",x"0099",x"007C",x"0013",
    x"0084",x"001B",x"00BB",x"0080",x"0312",x"00B5",x"00B5",x"0312",
    x"0080",x"0312",x"0052",x"003F",x"004C",x"004C",x"0084",x"00BB",
    x"0015",x"02A0",x"0080",x"0204",x"02FA",x"0268",x"0220",x"0006",
    x"02A1",x"0089",x"0204",x"02F3",x"03B9",x"000F",x"0271",x"0049",
    x"0001",x"02F9",x"00EC",x"0026",x"0288",x"0268",x"0009",x"0288",
    x"0268",x"02B8",x"0028",x"0268",x"02B1",x"0001",x"02F9",x"00F9",
    x"0040",x"028A",x"00AB",x"0004",x"01E8",x"0174",x"0013",x"02B8",
    x"0029",x"0258",x"0200",x"02D3",x"00AB",x"0004",x"017C",x"03AF",
    x"02B8",x"003D",x"0258",x"000B",x"0004",x"017C",x"0378",x"0200",
    x"02C6",x"00AB",x"0004",x"017C",x"03AF",x"0200",x"02C0",x"02A1",
    x"0089",x"0204",x"02BC",x"0275",x"02BA",x"000C",x"02B8",x"0006",
    x"0004",x"01EC",x"03E0",x"014A",x"020B",x"0006",x"0001",x"02BA",
    x"00BB",x"0026",x"0200",x"0007",x"0285",x"02F0",x"02FD",x"000C",
    x"0111",x"0001",x"02AA",x"0011",x"004D",x"00D1",x"02BA",x"0004",
    x"02B5",x"028B",x"026B",x"0009",x"0012",x"022C",x"0005",x"0200",
    x"0296",x"02A0",x"0268",x"0200",x"0292",x"00AB",x"0004",x"017C",
    x"0378",x"02A0",x"0080",x"0204",x"028A",x"0014",x"0014",x"0004",
    x"01E8",x"00C5",x"000C",x"02A0",x"0080",x"0204",x"0280",x"0014",
    x"02B8",x"002C",x"0258",x"000B",x"0220",x"000F",x"02A0",x"0268",
    x"02B8",x"003D",x"0268",x"00AB",x"0004",x"01E8",x"01A3",x"009D",
    x"02B8",x"0020",x"0268",x"02B8",x"0054",x"0268",x"02B8",x"004F",
    x"0268",x"02B8",x"0020",x"0268",x"00AB",x"0004",x"01E8",x"01A3",
    x"0200",x"025D",x"00AB",x"0004",x"01E8",x"016B",x"0200",x"0257",
    x"0015",x"02B8",x"0028",x"0268",x"00AB",x"0004",x"01E8",x"01A3",
    x"02A0",x"0004",x"01E8",x"0158",x"02FB",x"0002",x"0004",x"01E8",
    x"01A3",x"02B8",x"0029",x"0258",x"000B",x"0285",x"0354",x"02FD",
    x"002D",x"0275",x"00A9",x"0011",x"0289",x"0001",x"02F9",x"00AF",
    x"0040",x"02BA",x"0003",x"014C",x"0203",x"0005",x"02A0",x"0268",
    x"000A",x"0220",x"0007",x"037A",x"0003",x"0204",x"0227",x"01C0",
    x"0268",x"02B4",x"0014",x"0262",x"0220",x"011D",x"00AB",x"0014",
    x"0004",x"01E8",x"00C5",x"0200",x"021A",x"0275",x"0001",x"02BD",
    x"0078",x"0040",x"00A0",x"0268",x"0040",x"0268",x"0004",x"01E8",
    x"0229",x"0080",x"0204",x"0004",x"0378",x"000D",x"022C",x"0009",
    x"0274",x"0014",x"00A2",x"01C0",x"009D",x"0268",x"0001",x"037D",
    x"00AF",x"0040",x"022B",x"0006",x"00AB",x"0013",x"01E4",x"0001",
    x"037A",x"00B1",x"0040",x"0204",x"0046",x"0004",x"01E8",x"0265",
    x"0290",x"0378",x"0080",x"0204",x"0048",x"0378",x"00A3",x"0204",
    x"003A",x"0378",x"00B1",x"0204",x"0036",x"0378",x"00A4",x"0204",
    x"0032",x"0378",x"0001",x"0204",x"002E",x"0378",x"00A8",x"0204",
    x"002A",x"0378",x"000D",x"0204",x"0026",x"03B8",x"00E0",x"0378",
    x"0080",x"020C",x"002A",x"0290",x"0378",x"008A",x"020C",x"0007",
    x"0270",x"000C",x"0004",x"01E8",x"0158",x"0200",x"0036",x"0378",
    x"0084",x"020C",x"0002",x"0200",x"0030",x"0378",x"0082",x"020C",
    x"0010",x"0004",x"01E8",x"0158",x"0012",x"0004",x"01E8",x"0265",
    x"0004",x"01E8",x"023C",x"0004",x"01E8",x"02B4",x"00A3",x"02B4",
    x"02B7",x"0270",x"000C",x"0200",x"0018",x"0004",x"01E8",x"023C",
    x"00A4",x"0224",x"005B",x"02B0",x"0014",x"0378",x"008A",x"020C",
    x"0007",x"02B8",x"0084",x"0004",x"01E8",x"0158",x"0220",x"000F",
    x"0004",x"01E8",x"0158",x"0220",x"006D",x"0012",x"0220",x"0070",
    x"0275",x"0080",x"020C",x"0003",x"02B5",x"0200",x"0180",x"0085",
    x"03BD",x"001F",x"0015",x"0001",x"02FD",x"0096",x"002B",x"02A8",
    x"0258",x"0013",x"02B7",x"0275",x"0001",x"02A2",x"004A",x"0062",
    x"0004",x"01E8",x"0174",x"02B7",x"0275",x"0001",x"02B9",x"0010",
    x"0027",x"014A",x"0203",x"000A",x"0272",x"02BA",x"000A",x"0004",
    x"011C",x"01FB",x"02B2",x"0081",x"0220",x"000C",x"0088",x"0091",
    x"0082",x"0272",x"0004",x"011C",x"01FB",x"02F8",x"0030",x"0258",
    x"000B",x"02B0",x"0271",x"0081",x"02BA",x"000A",x"0004",x"011C",
    x"01FB",x"0081",x"02B2",x"0089",x"022C",x"0017",x"02B8",x"0020",
    x"0258",x"000B",x"02B7",x"0275",x"02A0",x"0080",x"020C",x"0003",
    x"02B5",x"0200",x"0134",x"0081",x"03B9",x"00C0",x"0379",x"00C0",
    x"020C",x"0040",x"0081",x"03B9",x"003F",x"02BA",x"0016",x"02B8",
    x"0004",x"0004",x"01EC",x"03E0",x"0151",x"0203",x"0007",x"0049",
    x"0001",x"02F9",x"00EC",x"0026",x"0200",x"0009",x"0111",x"0285",
    x"02F0",x"02FD",x"0008",x"0001",x"02A8",x"0049",x"00C1",x"0288",
    x"0258",x"000B",x"0009",x"0288",x"0258",x"000B",x"02B8",x"0028",
    x"0258",x"000B",x"02A0",x"0378",x"0080",x"0204",x"0006",x"0014",
    x"0200",x"000B",x"0270",x"0220",x"008F",x"0004",x"01E8",x"01FD",
    x"02B8",x"0029",x"0258",x"000B",x"02B7",x"02A0",x"0258",x"000B",
    x"0220",x"0009",x"0378",x"0080",x"020C",x"0004",x"0004",x"01E8",
    x"01FD",x"02B7",x"0258",x"000B",x"02B7",x"0275",x"0004",x"01EC",
    x"0049",x"02A0",x"0270",x"00A1",x"0282",x"035C",x"0004",x"01EC",
    x"0058",x"02B0",x"0082",x"0091",x"03BA",x"0007",x"0064",x"0064",
    x"03B9",x"0008",x"0204",x"0008",x"03B8",x"0003",x"02B9",x"0002",
    x"0110",x"0010",x"0200",x"0003",x"0110",x"0010",x"01C9",x"0274",
    x"009C",x"0004",x"0120",x"03EE",x"00A3",x"02B4",x"02FC",x"0004",
    x"02B7",x"0275",x"02A0",x"0378",x"0080",x"0204",x"0008",x"03B8",
    x"00C0",x"0378",x"00C0",x"0224",x"000A",x"0200",x"0002",x"02FC",
    x"0005",x"00A5",x"02A8",x"02B7",x"0275",x"0274",x"0094",x"0004",
    x"01E8",x"0229",x"01ED",x"0378",x"002D",x"020C",x"0001",x"000D",
    x"00A9",x"0272",x"0290",x"0378",x"0080",x"020C",x"0044",x"000A",
    x"0290",x"03B8",x"0008",x"0204",x"002B",x"02F9",x"0004",x"0290",
    x"0064",x"0064",x"03B8",x"0003",x"00C1",x"0290",x"03B8",x"0007",
    x"0204",x"0028",x"0009",x"0200",x"0025",x"0275",x"0274",x"0001",
    x"02BD",x"0078",x"0040",x"0001",x"02AC",x"00A1",x"0004",x"01E8",
    x"0229",x"0154",x"0204",x"0006",x"022B",x"0008",x"01C0",x"008A",
    x"02B4",x"02B7",x"0378",x"002D",x"022C",x"0010",x"0220",x"0008",
    x"0290",x"0064",x"0064",x"00C1",x"0290",x"03B8",x"0007",x"0204",
    x"0001",x"0009",x"000A",x"0290",x"03B8",x"0080",x"0204",x"000F",
    x"0009",x"0200",x"000C",x"03B8",x"00C0",x"0378",x"00C0",x"020C",
    x"0005",x"000A",x"02F9",x"0004",x"0220",x"0053",x"0009",x"02B2",
    x"0094",x"010B",x"0012",x"0272",x"0273",x"000B",x"00AD",x"0204",
    x"0004",x"02B8",x"002D",x"0258",x"000B",x"0004",x"01E8",x"01A3",
    x"02B3",x"02B2",x"02B4",x"02B7",x"0275",x"0284",x"0354",x"0001",
    x"037C",x"00AF",x"0040",x"0204",x"0020",x"02A0",x"0080",x"022C",
    x"0009",x"0014",x"00A5",x"02A9",x"0089",x"020C",x"0003",x"0008",
    x"0220",x"0006",x"00A5",x"00C5",x"02A8",x"0260",x"0001",x"037D",
    x"00AF",x"0040",x"022C",x"0007",x"00A5",x"01C0",x"0268",x"0001",
    x"037D",x"00AF",x"0040",x"022B",x"0006",x"02B7",x"02B5",x"0285",
    x"0354",x"00AA",x"02FA",x"0028",x"016A",x"0204",x"0004",x"02A8",
    x"0080",x"022C",x"0006",x"0015",x"02B8",x"000D",x"0268",x"02B7",
    x"0275",x"0272",x"0273",x"0004",x"01E8",x"030C",x"0272",x"0004",
    x"0174",x"01D4",x"02B1",x"02B5",x"02B8",x"0080",x"0268",x"0269",
    x"00AA",x"0281",x"035C",x"0275",x"0004",x"01EC",x"0058",x"02B3",
    x"02FB",x"0004",x"02B2",x"02B7",x"0275",x"0004",x"01EC",x"0049",
    x"0004",x"012C",x"03B7",x"0081",x"02B8",x"0007",x"0004",x"0114",
    x"02E6",x"015D",x"0275",x"0379",x"002D",x"0204",x"0006",x"0014",
    x"02B0",x"01C0",x"0270",x"0200",x"0005",x"0271",x"0004",x"01EC",
    x"00A5",x"02B1",x"0274",x"0004",x"01EC",x"003F",x"0224",x"0004",
    x"02B9",x"0006",x"0378",x"0045",x"020C",x"0002",x"02B9",x"0003",
    x"0001",x"02BA",x"00C5",x"0047",x"0251",x"01C9",x"008B",x"0013",
    x"02B4",x"0004",x"012C",x"03B7",x"0378",x"002E",x"0204",x"0036",
    x"0004",x"012C",x"01D2",x"0201",x"0039",x"0270",x"0001",x"02BD",
    x"00C5",x"0047",x"02A8",x"0141",x"020C",x"0003",x"02B0",x"0200",
    x"002D",x"02B0",x"0009",x"0271",x"0004",x"01EC",x"00A5",x"009B",
    x"020B",x"0001",x"000B",x"0273",x"0001",x"02BB",x"0005",x"0026",
    x"0004",x"01E0",x"00BB",x"0014",x"02A0",x"0338",x"0030",x"0001",
    x"02BB",x"00D4",x"0047",x"0004",x"01EC",x"0340",x"01C0",x"0004",
    x"01E0",x"0059",x"02B3",x"02B1",x"0220",x"003C",x"01DB",x"0271",
    x"0004",x"01EC",x"00A5",x"02B1",x"0220",x"0044",x"0014",x"0004",
    x"01EC",x"003F",x"0224",x"0004",x"0089",x"020C",x"0001",x"0009",
    x"004D",x"004D",x"009B",x"0203",x"0001",x"01DB",x"01D9",x"0378",
    x"0045",x"020C",x"0077",x"0274",x"0004",x"012C",x"03B7",x"0004",
    x"0170",x"008C",x"0221",x"0007",x"0004",x"012C",x"01D2",x"0209",
    x"0003",x"02B4",x"0200",x"0066",x"02B4",x"008A",x"0004",x"01EC",
    x"00A5",x"0004",x"012C",x"03B7",x"0004",x"0170",x"008C",x"0201",
    x"0003",x"0014",x"03FA",x"0040",x"03FA",x"0040",x"0272",x"0004",
    x"01EC",x"00A5",x"01DB",x"02A0",x"0004",x"012C",x"01D2",x"0221",
    x"0006",x"0338",x"0030",x"0082",x"0004",x"01EC",x"00A5",x"0098",
    x"02B9",x"000A",x"0093",x"0004",x"011C",x"01DC",x"00D3",x"02A0",
    x"0004",x"012C",x"01D2",x"0229",x"0013",x"02B2",x"037B",x"000A",
    x"020B",x"0002",x"03FA",x"0080",x"0272",x"03BA",x"0040",x"0204",
    x"0001",x"0023",x"02B1",x"008A",x"03F9",x"0008",x"03BA",x"0007",
    x"0271",x"0065",x"0065",x"03BA",x"0003",x"03B9",x"0003",x"009D",
    x"00CD",x"0115",x"0015",x"0113",x"037D",x"0048",x"020B",x"0005",
    x"033D",x"0048",x"012B",x"0200",x"000A",x"0001",x"037D",x"00BA",
    x"00FF",x"0203",x"0004",x"02FD",x"0046",x"0025",x"00EB",x"02B1",
    x"0200",x"0001",x"0023",x"0271",x"0014",x"0281",x"035C",x"008A",
    x"02FA",x"0015",x"0004",x"01EC",x"005C",x"0098",x"0004",x"01EC",
    x"006A",x"0001",x"02BB",x"00E2",x"0047",x"0004",x"01E0",x"00BB",
    x"02B1",x"008A",x"02B0",x"0080",x"0204",x"0006",x"0281",x"035C",
    x"0288",x"03F8",x"0080",x"0248",x"0004",x"01EC",x"003F",x"0223",
    x"0004",x"0014",x"0004",x"0324",x"014F",x"0034",x"0034",x"0275",
    x"01ED",x"0004",x"012C",x"03B7",x"0378",x"002E",x"0004",x"0378",
    x"023F",x"0275",x"0285",x"035C",x"02B8",x"0040",x"0268",x"01C0",
    x"0268",x"0001",x"037D",x"00D4",x"0047",x"022C",x"0006",x"02B7",
    x"02B8",x"0004",x"0200",x"0002",x"02B8",x"0007",x"0275",x"0274",
    x"008D",x"0094",x"00C2",x"02A8",x"0260",x"0154",x"022C",x"0004",
    x"02B4",x"02B7",x"0275",x"0081",x"0280",x"015D",x"03B8",x"00BF",
    x"0089",x"0203",x"0003",x"03F8",x"0040",x"0021",x"0240",x"015D",
    x"02B8",x"0001",x"0283",x"035C",x"0004",x"01EC",x"0340",x"01D2",
    x"0090",x"0004",x"0114",x"0345",x"0083",x"0188",x"0204",x"0017",
    x"0093",x"004F",x"004B",x"0113",x"0001",x"02FB",x"0005",x"0026",
    x"0285",x"015D",x"03BD",x"0040",x"0204",x"0002",x"02FB",x"0031",
    x"0271",x"0272",x"0004",x"01E0",x"00BB",x"02B2",x"02B1",x"000A",
    x"037A",x"0007",x"022C",x"0023",x"02B7",x"0275",x"02B8",x"0032",
    x"0004",x"017C",x"039A",x"02B7",x"0275",x"0001",x"02BA",x"0005",
    x"0023",x"0272",x"0004",x"0178",x"03AB",x"0089",x"020C",x"000B",
    x"0283",x"0163",x"02FB",x"0200",x"02B8",x"0010",x"0040",x"03D8",
    x"0258",x"02B0",x"02B7",x"0379",x"001F",x"020E",x"00C4",x"0379",
    x"000D",x"022E",x"0012",x"0204",x"00C4",x"0379",x"0008",x"0204",
    x"0085",x"0379",x"000C",x"0204",x"0167",x"0379",x"000A",x"0225",
    x"0020",x"0283",x"0163",x"02FB",x"0200",x"0004",x"01EC",x"0299",
    x"0280",x"0165",x"0080",x"0204",x"004E",x"009C",x"0282",x"0167",
    x"02FA",x"0200",x"0162",x"020E",x"0011",x"02B0",x"0270",x"0258",
    x"02B8",x"000D",x"0282",x"0165",x"0001",x"02FA",x"0085",x"0040",
    x"0250",x"000A",x"01C0",x"0250",x"0200",x"000D",x"02A0",x"02B5",
    x"0275",x"0168",x"022C",x"0019",x"009A",x"00A3",x"0284",x"0165",
    x"0004",x"01EC",x"02B1",x"0379",x"000A",x"020C",x"000F",x"033B",
    x"0200",x"0098",x"0008",x"0004",x"01EC",x"02E3",x"0283",x"0167",
    x"0153",x"020E",x"000A",x"009A",x"0200",x"0007",x"0280",x"0164",
    x"0338",x"0014",x"0004",x"01EC",x"02E3",x"0093",x"0243",x"0163",
    x"0280",x"015D",x"03B8",x"00EF",x"0240",x"015D",x"01C0",x"0240",
    x"0165",x"0200",x"001F",x"033B",x"0214",x"0379",x"000B",x"0204",
    x"0002",x"02FB",x"0028",x"0280",x"0166",x"0143",x"020D",x"0001",
    x"0083",x"0098",x"0004",x"01EC",x"02E3",x"02FA",x"0028",x"0153",
    x"0206",x"0002",x"033B",x"0014",x"0280",x"0167",x"0143",x"0206",
    x"0001",x"0083",x"02FB",x"0200",x"0200",x"011F",x"0280",x"0163",
    x"0004",x"01EC",x"02E3",x"0283",x"0163",x"015A",x"0224",x"00A7",
    x"02FB",x"0200",x"0004",x"01EC",x"0299",x"0013",x"0280",x"0166",
    x"02F8",x"0200",x"0143",x"020D",x"0001",x"000B",x"0281",x"0165",
    x"0089",x"0204",x"0016",x"0200",x"0006",x"0280",x"015D",x"03B8",
    x"00EF",x"0240",x"015D",x"02B8",x"0020",x"0011",x"0241",x"0165",
    x"0001",x"02F9",x"0086",x"0040",x"0248",x"02B8",x"0022",x"0040",
    x"0258",x"0200",x"00EA",x"0280",x"0165",x"0378",x"0027",x"022D",
    x"00D8",x"0283",x"0163",x"02FB",x"0200",x"0004",x"01EC",x"0299",
    x"0379",x"0060",x"0205",x"0002",x"0339",x"0020",x"0283",x"0163",
    x"0282",x"0167",x"0153",x"020C",x"000F",x"0004",x"0178",x"03C7",
    x"0283",x"0163",x"033B",x"0014",x"0243",x"0163",x"0280",x"0164",
    x"0338",x"0014",x"0240",x"0164",x"0280",x"0165",x"0080",x"020C",
    x"0022",x"008C",x"0098",x"0004",x"01EC",x"02E3",x"0153",x"020D",
    x"000C",x"0273",x"0004",x"01EC",x"030F",x"02B3",x"02FB",x"0200",
    x"02B0",x"0270",x"0258",x"033B",x"0200",x"00A1",x"0242",x"0164",
    x"0153",x"0204",x"0008",x"01E4",x"02FA",x"0200",x"02FB",x"0200",
    x"0004",x"01EC",x"02B1",x"0284",x"0165",x"000C",x"0244",x"0165",
    x"0001",x"02FC",x"0084",x"0040",x"0261",x"0283",x"0163",x"02FB",
    x"0200",x"0298",x"0379",x"000D",x"0204",x"0012",x"0339",x"0020",
    x"004D",x"0049",x"0041",x"03F9",x"0022",x"0041",x"0259",x"000B",
    x"02B5",x"0275",x"0168",x"020C",x"0001",x"0258",x"0200",x"0075",
    x"01C0",x"0260",x"02B0",x"0270",x"0258",x"033B",x"0200",x"0098",
    x"0004",x"01EC",x"02E3",x"0280",x"0166",x"0142",x"020C",x"000F",
    x"02FA",x"0200",x"0290",x"02B5",x"0275",x"0168",x"020C",x"0003",
    x"02B0",x"0270",x"0250",x"033A",x"0200",x"02FA",x"0014",x"0242",
    x"0163",x"02FB",x"0200",x"02FA",x"0200",x"009D",x"000D",x"02B8",
    x"0022",x"0040",x"0155",x"0204",x"0003",x"0268",x"0220",x"0005",
    x"0280",x"015D",x"03B8",x"00EF",x"0240",x"015D",x"01C0",x"0240",
    x"0165",x"0093",x"0200",x"0039",x"0281",x"0165",x"0379",x"0027",
    x"022D",x"0189",x"0283",x"0163",x"0281",x"0167",x"014B",x"0205",
    x"000D",x"0004",x"0178",x"03C7",x"0280",x"0164",x"0338",x"0014",
    x"0240",x"0164",x"0283",x"0163",x"033B",x"0014",x"02FB",x"0200",
    x"0004",x"01EC",x"0299",x"000B",x"0284",x"0165",x"00A4",x"0204",
    x"0014",x"0013",x"0298",x"02B5",x"0275",x"0168",x"020C",x"0007",
    x"000B",x"0258",x"0013",x"02B8",x"0022",x"0040",x"0258",x"000B",
    x"009A",x"0012",x"0004",x"01EC",x"02B1",x"0004",x"01EC",x"027E",
    x"033B",x"0200",x"0243",x"0163",x"02B0",x"02B7",x"0275",x"0285",
    x"0162",x"03BD",x"0001",x"0298",x"0001",x"0378",x"0005",x"0023",
    x"0204",x"0005",x"0040",x"03B8",x"0010",x"0200",x"0006",x"02B8",
    x"0022",x"0040",x"0258",x"02B8",x"0020",x"01C5",x"0245",x"0162",
    x"02B7",x"0275",x"029D",x"0001",x"03BD",x"00FF",x"002F",x"0280",
    x"0162",x"03B8",x"0030",x"0378",x"0020",x"0204",x"0004",x"0040",
    x"01E8",x"0200",x"0004",x"0001",x"02B8",x"0005",x"0023",x"0258",
    x"02B7",x"0275",x"0280",x"0354",x"0270",x"00C4",x"0095",x"02A8",
    x"0001",x"0378",x"0005",x"0023",x"020C",x"0004",x"02B8",x"000D",
    x"0200",x"0015",x"0064",x"0060",x"03B8",x"003F",x"0082",x"02F8",
    x"0020",x"004E",x"004A",x"0042",x"03FA",x"0022",x"0042",x"0015",
    x"026A",x"0001",x"037C",x"00AC",x"0040",x"0203",x"0001",x"0260",
    x"015D",x"0225",x"0023",x"01C0",x"0260",x"0014",x"02B0",x"0104",
    x"0244",x"0165",x"02B7",x"0275",x"0282",x"0166",x"0150",x"020E",
    x"0002",x"01C9",x"02B7",x"0081",x"02F9",x"0200",x"02FA",x"0200",
    x"0288",x"0001",x"03F8",x"0005",x"0023",x"0001",x"03B8",x"00FF",
    x"000F",x"0204",x"0007",x"0011",x"0151",x"022D",x"000E",x"033A",
    x"0200",x"02B7",x"0339",x"0200",x"02BA",x"0014",x"0004",x"011C",
    x"01FB",x"0008",x"004C",x"0082",x"004E",x"00C2",x"02B7",x"0275",
    x"0273",x"02FB",x"0200",x"0282",x"0166",x"02FA",x"0200",x"0298",
    x"0001",x"0378",x"0005",x"0023",x"0204",x"0004",x"0013",x"015A",
    x"0225",x"000A",x"02B8",x"0022",x"0040",x"0258",x"02B3",x"0098",
    x"0004",x"03EC",x"02E4",x"0275",x"02BD",x"0162",x"02B8",x"0020",
    x"0268",x"004C",x"004C",x"0268",x"01C0",x"0268",x"0268",x"0268",
    x"02B8",x"00DC",x"0268",x"02B8",x"0078",x"0240",x"00F8",x"02B7",
    x"0275",x"0080",x"0204",x"0024",x"02BD",x"0004",x"0082",x"0090",
    x"0040",x"03B8",x"00F0",x"020C",x"0005",x"0015",x"004E",x"004E",
    x"0220",x"000A",x"03FD",x"0040",x"025D",x"009D",x"000D",x"0042",
    x"026A",x"0042",x"026A",x"01D2",x"026A",x"0282",x"015D",x"03BA",
    x"0080",x"0204",x"0004",x"01D2",x"026A",x"026A",x"026A",x"02B7",
    x"009D",x"02B8",x"0040",x"0268",x"01C0",x"0268",x"0268",x"0268",
    x"0220",x"0014",x"0275",x"0273",x"0001",x"02BC",x"0065",x"0047",
    x"0274",x"02B8",x"0010",x"0004",x"0114",x"0338",x"02BB",x"000C",
    x"02BA",x"0002",x"0004",x"01E4",x"037D",x"02B4",x"02B9",x"0040",
    x"0378",x"0002",x"0204",x"0002",x"02B9",x"0080",x"0261",x"02B9",
    x"0018",x"0261",x"02B3",x"0263",x"0043",x"0263",x"000C",x"02B9",
    x"0050",x"0261",x"000C",x"0261",x"033C",x"0008",x"02B7",x"0275",
    x"02B8",x"000C",x"0004",x"01EC",x"03E0",x"00A4",x"020C",x"0009",
    x"0001",x"02BC",x"000B",x"0041",x"0001",x"02A0",x"000C",x"0080",
    x"02B7",x"0014",x"02A0",x"00C4",x"033C",x"0003",x"0220",x"000B",
    x"0275",x"0283",x"0163",x"02FB",x"0200",x"0004",x"01EC",x"0299",
    x"0283",x"0166",x"0243",x"0163",x"02FB",x"0200",x"0004",x"01EC",
    x"027E",x"02B7",x"0275",x"0274",x"02B8",x"0008",x"0004",x"0114",
    x"0338",x"033C",x"0004",x"0261",x"0274",x"02BB",x"0034",x"02BA",
    x"007F",x"0004",x"01E4",x"037D",x"02B4",x"0260",x"02B3",x"02B7",
    x"0275",x"0274",x"0034",x"0273",x"0272",x"0271",x"0034",x"0001",
    x"02BB",x"0001",x"00C0",x"0270",x"0004",x"0120",x"001F",x"02B0",
    x"02A1",x"0379",x"01C1",x"020C",x"0003",x"0004",x"01C0",x"0040",
    x"02B1",x"0034",x"02B2",x"02B3",x"02B4",x"0034",x"02B7",x"00E1");

  CONSTANT INIT_VOICE : arr8 := (
    x"E8",x"BB",x"E8",x"87",x"E8",x"17",x"E8",x"37",x"E8",x"F7",x"E8",x"8F",x"E8",x"CF",x"E2",x"D8",
    x"E2",x"9A",x"E2",x"89",x"E2",x"DD",x"E2",x"37",x"E2",x"2F",x"EA",x"04",x"EA",x"54",x"EA",x"4C",
    x"EA",x"D2",x"EA",x"8A",x"EA",x"8E",x"EA",x"B1",x"EA",x"FD",x"EA",x"53",x"EA",x"AB",x"EA",x"47",
    x"EA",x"CF",x"EA",x"FF",x"E6",x"10",x"E6",x"48",x"E6",x"3C",x"E6",x"62",x"E6",x"8A",x"E6",x"BA",
    x"E6",x"76",x"E6",x"5E",x"E6",x"C1",x"E6",x"B1",x"E6",x"CB",x"EE",x"C8",x"EE",x"98",x"EE",x"F8",
    x"EE",x"C2",x"EE",x"1E",x"EE",x"7E",x"EE",x"2D",x"EE",x"6D",x"EE",x"1D",x"EE",x"5D",x"EE",x"3D",
    x"18",x"2B",x"15",x"C0",x"39",x"24",x"43",x"E2",x"1F",x"00",x"18",x"23",x"24",x"C0",x"28",x"23",
    x"62",x"C6",x"1D",x"A5",x"03",x"20",x"66",x"52",x"0C",x"95",x"03",x"00",x"19",x"2C",x"0C",x"80",
    x"31",x"12",x"62",x"A7",x"1C",x"00",x"18",x"2C",x"0C",x"C0",x"29",x"94",x"E0",x"64",x"9C",x"85",
    x"02",x"38",x"85",x"12",x"9C",x"8C",x"03",x"00",x"10",x"35",x"E7",x"55",x"AD",x"6D",x"7F",x"26",
    x"91",x"85",x"D4",x"3C",x"AB",x"D6",x"CF",x"99",x"7A",x"00",x"10",x"34",x"6F",x"A1",x"86",x"CF",
    x"3E",x"AB",x"0D",x"BB",x"86",x"7C",x"6C",x"B5",x"6D",x"CF",x"24",x"B2",x"88",x"9E",x"A7",x"16",
    x"F3",x"A9",x"D2",x"E6",x"3D",x"D5",x"55",x"FD",x"01",x"00",x"10",x"32",x"74",x"98",x"A9",x"B7",
    x"81",x"1E",x"A9",x"87",x"F4",x"66",x"A3",x"FC",x"8B",x"D2",x"96",x"94",x"FB",x"FF",x"10",x"03",
    x"80",x"8E",x"16",x"0D",x"00",x"10",x"32",x"7C",x"90",x"AB",x"B7",x"81",x"1E",x"A9",x"A7",x"6E",
    x"F7",x"22",x"DD",x"C7",x"AA",x"FE",x"A5",x"9C",x"DE",x"CC",x"7E",x"F4",x"2E",x"AC",x"FA",x"C7",
    x"D9",x"91",x"A5",x"A5",x"E4",x"DC",x"5F",x"F4",x"2B",x"9D",x"FC",x"03",x"00",x"10",x"31",x"8F",
    x"DC",x"FF",x"8C",x"7C",x"97",x"F6",x"41",x"E6",x"E3",x"F4",x"F4",x"F6",x"47",x"23",x"C2",x"84",
    x"B6",x"85",x"74",x"FF",x"D0",x"DD",x"CF",x"EE",x"3F",x"B7",x"EB",x"01",x"00",x"74",x"7B",x"A3",
    x"DC",x"2D",x"3A",x"5A",x"B7",x"56",x"EE",x"45",x"DF",x"5B",x"DA",x"BF",x"68",x"E9",x"3B",x"FD",
    x"1F",x"F5",x"78",x"27",x"FF",x"A2",x"4E",x"F2",x"DC",x"1F",x"00",x"10",x"36",x"76",x"9B",x"A9",
    x"B7",x"BD",x"1A",x"1F",x"66",x"D4",x"85",x"A3",x"BB",x"CB",x"95",x"83",x"00",x"10",x"32",x"6E",
    x"DA",x"27",x"BB",x"7D",x"22",x"1F",x"C6",x"94",x"16",x"9C",x"DE",x"97",x"D6",x"A5",x"D3",x"7F",
    x"52",x"72",x"58",x"F2",x"4F",x"D7",x"85",x"03",x"00",x"10",x"32",x"35",x"96",x"A9",x"B9",x"BD",
    x"1A",x"1F",x"86",x"CE",x"6E",x"13",x"3D",x"09",x"E9",x"F6",x"00",x"10",x"32",x"7B",x"94",x"AB",
    x"B7",x"81",x"1E",x"A9",x"87",x"6E",x"AF",x"1B",x"DD",x"F9",x"AA",x"FE",x"A4",x"57",x"E6",x"CC",
    x"5E",x"F4",x"36",x"AD",x"FA",x"C7",x"D5",x"B5",x"A4",x"A5",x"ED",x"DC",x"5F",x"F4",x"73",x"9E",
    x"FC",x"03",x"00",x"10",x"32",x"F7",x"9F",x"A9",x"BD",x"3F",x"22",x"11",x"86",x"6E",x"CF",x"A3",
    x"DB",x"FB",x"46",x"EB",x"C8",x"E9",x"3F",x"00",x"10",x"32",x"AC",x"98",x"27",x"BD",x"81",x"22",
    x"1F",x"87",x"AE",x"7E",x"1C",x"6D",x"81",x"E7",x"FF",x"72",x"E4",x"20",x"00",x"F1",x"E1",x"00",
    x"00",x"11",x"FC",x"13",x"FF",x"13",x"FF",x"00",x"FE",x"13",x"FF",x"00",x"11",x"FF",x"00",x"FF",
    x"00",x"F7",x"00",x"18",x"32",x"DD",x"A0",x"7D",x"81",x"0F",x"C7",x"03",x"E3",x"EA",x"53",x"C6",
    x"75",x"AB",x"F0",x"41",x"E8",x"9E",x"17",x"73",x"A1",x"D2",x"DC",x"62",x"F6",x"14",x"34",x"4D",
    x"0F",x"8C",x"B7",x"54",x"99",x"5A",x"CB",x"5F",x"80",x"84",x"6D",x"88",x"F3",x"65",x"2A",x"73",
    x"BD",x"F5",x"77",x"50",x"AD",x"5D",x"EF",x"A1",x"5A",x"F5",x"45",x"3C",x"80",x"53",x"14",x"83",
    x"C8",x"BC",x"C9",x"05",x"60",x"09",x"03",x"68",x"B0",x"AF",x"A9",x"81",x"00",x"38",x"78",x"D8",
    x"8F",x"D9",x"61",x"A2",x"35",x"77",x"90",x"7F",x"07",x"D3",x"DA",x"80",x"FF",x"EC",x"B4",x"66",
    x"DF",x"31",x"D8",x"D8",x"89",x"BF",x"65",x"9B",x"9D",x"5E",x"82",x"3E",x"12",x"24",x"21",x"6F",
    x"FC",x"24",x"83",x"03",x"00",x"F2",x"F3",x"1F",x"5C",x"3E",x"48",x"90",x"60",x"0D",x"EE",x"03",
    x"A5",x"8B",x"00",x"00",x"1A",x"FD",x"38",x"50",x"A6",x"00",x"F0",x"03",x"21",x"6E",x"C7",x"8D",
    x"D9",x"F3",x"A0",x"30",x"D2",x"6F",x"22",x"F1",x"1A",x"95",x"71",x"89",x"0C",x"44",x"8A",x"C6",
    x"A7",x"D1",x"6B",x"A2",x"33",x"AF",x"9A",x"41",x"D1",x"CE",x"FC",x"2E",x"3B",x"4D",x"74",x"C6",
    x"24",x"13",x"18",x"91",x"61",x"9E",x"94",x"D7",x"75",x"CE",x"D4",x"53",x"0A",x"24",x"2A",x"DB",
    x"8F",x"F2",x"34",x"D0",x"19",x"5B",x"6A",x"80",x"64",x"47",x"79",x"D7",x"2D",x"F7",x"39",x"53",
    x"4B",x"09",x"90",x"C8",x"68",x"1F",x"AB",x"BD",x"46",x"69",x"DA",x"26",x"85",x"08",x"A2",x"FE",
    x"71",x"F1",x"55",x"A9",x"A4",x"74",x"E0",x"87",x"0F",x"1E",x"65",x"CC",x"DC",x"48",x"06",x"2C",
    x"2A",x"F3",x"DB",x"E6",x"B8",x"52",x"9A",x"7D",x"A8",x"A0",x"46",x"85",x"7E",x"97",x"0D",x"47",
    x"3A",x"63",x"FB",x"D4",x"2B",x"B0",x"28",x"BE",x"50",x"C2",x"44",x"67",x"DE",x"A1",x"88",x"16",
    x"19",x"E6",x"53",x"39",x"96",x"28",x"3F",x"86",x"49",x"05",x"80",x"C7",x"06",x"10",x"49",x"27",
    x"71",x"00",x"10",x"C9",x"F8",x"46",x"DB",x"33",x"5F",x"51",x"FB",x"00",x"0B",x"CE",x"76",x"9F",
    x"68",x"36",x"A6",x"0D",x"B2",x"67",x"A8",x"59",x"19",x"A6",x"0A",x"D8",x"57",x"2A",x"30",x"84",
    x"24",x"E0",x"22",x"32",x"8D",x"6B",x"B4",x"CF",x"60",x"B3",x"F4",x"DF",x"DF",x"82",x"C5",x"A0",
    x"69",x"91",x"0C",x"7A",x"76",x"AC",x"1F",x"C9",x"42",x"AD",x"32",x"AF",x"98",x"41",x"8B",x"8A",
    x"F5",x"37",x"59",x"8A",x"75",x"C6",x"DE",x"63",x"C8",x"D8",x"C9",x"1E",x"57",x"C3",x"91",x"CE",
    x"B8",x"88",x"EE",x"15",x"22",x"8B",x"13",x"0E",x"B3",x"D0",x"7D",x"68",x"03",x"F3",x"FB",x"18",
    x"23",x"1C",x"00",x"29",x"18",x"80",x"2A",x"B9",x"A6",x"2E",x"22",x"20",x"D9",x"C1",x"1D",x"36",
    x"63",x"99",x"CE",x"D4",x"46",x"04",x"22",x"33",x"BA",x"C7",x"6A",x"B6",x"CE",x"C9",x"EF",x"D7",
    x"0B",x"24",x"58",x"44",x"A7",x"A1",x"9D",x"FA",x"4D",x"44",x"12",x"47",x"20",x"5D",x"9C",x"32",
    x"2F",x"54",x"C9",x"0A",x"13",x"FA",x"27",x"3C",x"E9",x"34",x"E4",x"02",x"B0",x"26",x"52",x"40",
    x"98",x"93",x"58",x"00",x"C5",x"64",x"8E",x"86",x"7B",x"91",x"07",x"00",x"93",x"38",x"D0",x"F1",
    x"1F",x"E2",x"01",x"58",x"F3",x"39",x"70",x"9E",x"6B",x"EC",x"9E",x"80",x"92",x"1D",x"FE",x"6D",
    x"F5",x"9C",x"67",x"65",x"09",x"E0",x"00",x"00",x"00",x"F1",x"D0",x"DC",x"3C",x"06",x"1C",x"4C",
    x"6E",x"07",x"FC",x"B1",x"54",x"9A",x"DA",x"A7",x"60",x"41",x"A4",x"EB",x"7D",x"A1",x"95",x"2A",
    x"C3",x"16",x"11",x"14",x"D0",x"6C",x"0D",x"1F",x"A6",x"50",x"6B",x"38",x"27",x"82",x"82",x"99",
    x"9D",x"FF",x"C7",x"1C",x"A3",x"4C",x"97",x"34",x"50",x"53",x"95",x"00",x"AA",x"E6",x"91",x"2D",
    x"19",x"00",x"10",x"F2",x"04",x"2F",x"DB",x"D0",x"06",x"F1",x"00",x"10",x"33",x"66",x"A6",x"67",
    x"79",x"85",x"22",x"A9",x"87",x"E6",x"55",x"B5",x"6E",x"00",x"50",x"24",x"F5",x"CC",x"BC",x"67",
    x"9E",x"ED",x"0D",x"8A",x"A4",x"9E",x"51",x"9B",x"6B",x"F6",x"5F",x"BA",x"97",x"D1",x"EE",x"45",
    x"CF",x"BF",x"B9",x"3B",x"04",x"8D",x"39",x"F9",x"F9",x"7C",x"AE",x"48",x"EA",x"11",x"7D",x"7B",
    x"69",x"EE",x"A5",x"A6",x"31",x"BD",x"3F",x"1E",x"00",x"10",x"33",x"56",x"22",x"47",x"4D",x"81",
    x"AE",x"92",x"58",x"C6",x"85",x"53",x"68",x"D1",x"6F",x"95",x"EE",x"D7",x"D8",x"67",x"1C",x"35",
    x"F4",x"CE",x"12",x"F2",x"9A",x"FB",x"8D",x"D8",x"98",x"20",x"11",x"86",x"22",x"7A",x"3F",x"5E",
    x"FD",x"47",x"5B",x"57",x"BB",x"FF",x"28",x"4B",x"6B",x"F9",x"1F",x"2D",x"8F",x"ED",x"FE",x"F1",
    x"00",x"D0",x"56",x"10",x"33",x"EE",x"D4",x"E5",x"F9",x"BF",x"23",x"2D",x"67",x"B4",x"D5",x"92",
    x"DB",x"97",x"B6",x"68",x"52",x"FB",x"D1",x"F2",x"4F",x"62",x"4F",x"FA",x"71",x"CA",x"EB",x"47",
    x"39",x"5F",x"69",x"FD",x"E8",x"83",x"2D",x"AB",x"8F",x"07",x"00",x"D0",x"3E",x"18",x"33",x"ED",
    x"5E",x"F9",x"82",x"8A",x"D2",x"03",x"03",x"EB",x"14",x"C2",x"A6",x"5D",x"33",x"B5",x"26",x"D7",
    x"E2",x"C2",x"90",x"D6",x"86",x"B4",x"FB",x"D1",x"96",x"76",x"FA",x"4F",x"67",x"3A",x"63",x"C8",
    x"90",x"DA",x"F6",x"1E",x"35",x"B2",x"07",x"90",x"AF",x"CC",x"78",x"00",x"D0",x"61",x"D0",x"19",
    x"D0",x"55",x"F1",x"00",x"D0",x"61",x"10",x"37",x"76",x"99",x"AD",x"B3",x"7F",x"1E",x"A2",x"A7",
    x"74",x"8F",x"B3",x"1A",x"CC",x"ED",x"8D",x"A4",x"37",x"A8",x"DD",x"9F",x"EE",x"9E",x"1D",x"75",
    x"71",x"29",x"F7",x"A2",x"66",x"30",x"DD",x"7E",x"E5",x"00",x"98",x"23",x"C2",x"C7",x"03",x"00",
    x"D0",x"06",x"D0",x"06",x"D0",x"53",x"D0",x"06",x"F1",x"00",x"D0",x"06",x"D0",x"06",x"D0",x"A7",
    x"F1",x"00",x"10",x"32",x"F6",x"9F",x"A9",x"BD",x"3F",x"22",x"11",x"86",x"6E",x"CF",x"A3",x"BB",
    x"FB",x"46",x"EB",x"C8",x"E9",x"FF",x"3D",x"B4",x"15",x"F1",x"00",x"D8",x"B0",x"D8",x"B4",x"F1",
    x"00",x"D0",x"56",x"10",x"34",x"76",x"9B",x"AB",x"B9",x"BD",x"15",x"1F",x"87",x"EE",x"C6",x"1B",
    x"B5",x"3B",x"EB",x"FE",x"A3",x"A5",x"ED",x"DC",x"9F",x"8E",x"BC",x"9D",x"EB",x"96",x"E3",x"01",
    x"00",x"10",x"32",x"6D",x"A0",x"A7",x"BF",x"81",x"15",x"1F",x"CA",x"B4",x"B6",x"9B",x"1E",x"88",
    x"96",x"7D",x"53",x"FF",x"D3",x"77",x"8E",x"6A",x"00",x"7D",x"0A",x"F1",x"00",x"D0",x"56",x"10",
    x"32",x"9C",x"A0",x"A9",x"2D",x"BF",x"22",x"1F",x"68",x"F4",x"F4",x"A3",x"F8",x"93",x"DE",x"80",
    x"55",x"7F",x"D3",x"DA",x"AF",x"E6",x"4F",x"4A",x"03",x"56",x"1C",x"4A",x"CD",x"3C",x"7A",x"43",
    x"9C",x"99",x"77",x"4A",x"F9",x"CD",x"0B",x"4A",x"06",x"00",x"53",x"26",x"78",x"3C",x"00",x"D0",
    x"3E",x"D8",x"D2",x"FE",x"D0",x"56",x"D8",x"BA",x"F1",x"00",x"D0",x"61",x"D0",x"55",x"F3",x"D0",
    x"56",x"D8",x"BA",x"F1",x"00",x"D0",x"61",x"D8",x"9E",x"D0",x"61",x"F5",x"D0",x"56",x"D8",x"BA",
    x"F1",x"00",x"D0",x"06",x"D0",x"06",x"D0",x"53",x"D0",x"06",x"D0",x"06",x"F4",x"D0",x"56",x"D8",
    x"BA",x"F1",x"00",x"D0",x"06",x"D0",x"06",x"D8",x"D1",x"D0",x"56",x"D8",x"BA",x"F1",x"00",x"D8",
    x"CD",x"FE",x"D0",x"56",x"D8",x"BA",x"F1",x"00",x"D8",x"B0",x"D8",x"B4",x"D0",x"56",x"D8",x"BA",
    x"F1",x"00",x"D0",x"56",x"10",x"32",x"6D",x"93",x"AB",x"B1",x"BF",x"1A",x"1F",x"46",x"EE",x"ED",
    x"1A",x"AD",x"C7",x"6A",x"F6",x"A2",x"35",x"5B",x"DD",x"9F",x"F4",x"A4",x"9B",x"FC",x"DB",x"8B",
    x"3C",x"00",x"87",x"60",x"F6",x"7A",x"68",x"2B",x"D8",x"13",x"F1",x"00",x"D0",x"3E",x"D8",x"D2",
    x"D0",x"56",x"D8",x"13",x"F1",x"00",x"D0",x"61",x"D0",x"55",x"F3",x"D0",x"56",x"D8",x"13",x"F1",
    x"00",x"D0",x"61",x"D8",x"9E",x"D0",x"61",x"D0",x"56",x"D8",x"13",x"F1",x"00",x"D0",x"06",x"D0",
    x"06",x"D0",x"53",x"D0",x"06",x"D0",x"06",x"F4",x"D0",x"56",x"D8",x"13",x"F1",x"00",x"D0",x"06",
    x"D0",x"06",x"D8",x"D1",x"D0",x"56",x"D8",x"13",x"F1",x"00",x"D8",x"CD",x"F7",x"D0",x"56",x"D8",
    x"13",x"F1",x"00",x"D8",x"B0",x"D8",x"B4",x"D0",x"56",x"D8",x"13",x"F1",x"00",x"10",x"25",x"02",
    x"C0",x"10",x"97",x"BC",x"A4",x"01",x"A8",x"02",x"93",x"CF",x"D8",x"7D",x"B6",x"D6",x"FE",x"6A",
    x"7C",x"1C",x"D2",x"1D",x"D0",x"EE",x"3F",x"5A",x"FE",x"4D",x"FD",x"47",x"4B",x"C6",x"B9",x"FF",
    x"88",x"03",x"20",x"43",x"27",x"97",x"E9",x"40",x"3D",x"BD",x"ED",x"D5",x"F8",x"38",x"A3",x"2E",
    x"24",x"DD",x"5D",x"F4",x"CD",x"A4",x"DB",x"8F",x"BA",x"95",x"74",x"FF",x"D1",x"8E",x"72",x"EE",
    x"1F",x"0F",x"00",x"D0",x"3E",x"10",x"35",x"37",x"9A",x"AB",x"B5",x"BF",x"1A",x"1F",x"C7",x"74",
    x"4F",x"B3",x"FA",x"97",x"BE",x"7E",x"15",x"03",x"52",x"33",x"93",x"66",x"60",x"52",x"00",x"AC",
    x"F1",x"06",x"4E",x"1A",x"80",x"3B",x"06",x"C5",x"0C",x"F7",x"EA",x"69",x"ED",x"AF",x"C6",x"C7",
    x"21",x"ED",x"90",x"E7",x"06",x"A2",x"15",x"F6",x"D4",x"7F",x"3E",x"A4",x"00",x"48",x"E3",x"91",
    x"C7",x"03",x"00",x"D0",x"56",x"D8",x"BA",x"F1",x"00",x"D0",x"56",x"D8",x"13",x"F1",x"00",x"10",
    x"28",x"1D",x"C0",x"18",x"1D",x"7C",x"86",x"DC",x"33",x"B5",x"2E",x"4F",x"E3",x"D2",x"8C",x"D6",
    x"7F",x"75",x"F7",x"51",x"1B",x"B1",x"6E",x"3F",x"7A",x"FB",x"D5",x"FD",x"A1",x"0D",x"00",x"D0",
    x"06",x"F1",x"00",x"10",x"34",x"76",x"9C",x"A9",x"BB",x"7F",x"1D",x"22",x"68",x"74",x"7F",x"AB",
    x"FC",x"8F",x"B2",x"77",x"73",x"FF",x"99",x"CB",x"30",x"62",x"C7",x"5F",x"53",x"82",x"9E",x"4F",
    x"E2",x"01",x"58",x"F2",x"F1",x"67",x"4C",x"44",x"53",x"6F",x"FB",x"3A",x"44",x"90",x"A8",x"E9",
    x"4B",x"77",x"97",x"2B",x"D1",x"E3",x"01",x"00",x"D0",x"19",x"D0",x"55",x"F1",x"00",x"10",x"32",
    x"B4",x"A9",x"A9",x"BB",x"7F",x"1D",x"22",x"48",x"EE",x"96",x"0D",x"DD",x"8F",x"6B",x"FF",x"72",
    x"BB",x"73",x"E8",x"1E",x"6D",x"F9",x"17",x"7D",x"69",x"EB",x"FE",x"A1",x"2C",x"E3",x"DC",x"60",
    x"F4",x"B4",x"9B",x"1A",x"C4",x"9D",x"69",x"73",x"56",x"9B",x"A8",x"4B",x"45",x"37",x"88",x"63",
    x"AB",x"E2",x"01",x"00",x"F1",x"00",x"F1",x"00",x"F1",x"00",x"F1",x"00",x"F1",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00");

END PACKAGE;