library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity patrons_list is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0);
	lines : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of patrons_list is
	type rom is array(0 to  2519) of std_logic_vector(7 downto 0);
	signal rom_data: rom :=
	( --   0     1     2     3     4     5     6     7     8     9    10    11    12    13    14    15    16    17    18    19    20    21    22    23    24    25    26    27    28    29    30    31    32    33    34    35    36    37    38    39
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 0
		X"20",X"20",X"53",X"75",X"70",X"70",X"6F",X"72",X"74",X"20",X"61",X"74",X"20",X"68",X"74",X"74",X"70",X"73",X"3A",X"2F",X"2F",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 1
		X"20",X"20",X"63",X"61",X"74",X"61",X"72",X"73",X"65",X"2E",X"6D",X"65",X"2F",X"6D",X"75",X"6C",X"74",X"69",X"63",X"6F",X"72",X"65",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 2
		X"20",X"20",X"6F",X"72",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 3
		X"20",X"20",X"53",X"75",X"70",X"70",X"6F",X"72",X"74",X"20",X"61",X"74",X"20",X"68",X"74",X"74",X"70",X"73",X"3A",X"2F",X"2F",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 4
		X"20",X"20",X"77",X"77",X"77",X"2E",X"70",X"61",X"74",X"72",X"65",X"6F",X"6E",X"2E",X"63",X"6F",X"6D",X"2F",X"76",X"74",X"72",X"75",X"63",X"63",X"6F",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 5
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 6
		X"20",X"20",X"54",X"68",X"61",X"6E",X"6B",X"73",X"20",X"74",X"6F",X"20",X"6D",X"79",X"20",X"70",X"61",X"74",X"72",X"6F",X"6E",X"73",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 7
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 8
		X"20",X"20",X"41",X"6C",X"65",X"6E",X"63",X"61",X"72",X"20",X"53",X"75",X"63",X"65",X"6E",X"61",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 9
		X"20",X"20",X"41",X"6C",X"65",X"78",X"61",X"6E",X"64",X"72",X"65",X"20",X"47",X"75",X"69",X"6D",X"61",X"72",X"61",X"65",X"73",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 10
		X"20",X"20",X"41",X"6C",X"66",X"72",X"65",X"64",X"6F",X"20",X"4A",X"75",X"6E",X"69",X"6F",X"72",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 11
		X"20",X"20",X"41",X"6E",X"64",X"79",X"20",X"4D",X"63",X"43",X"61",X"6C",X"6C",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 12
		X"20",X"20",X"41",X"6E",X"64",X"79",X"20",X"50",X"61",X"6C",X"6D",X"65",X"72",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 13
		X"20",X"20",X"41",X"6E",X"74",X"6F",X"6E",X"69",X"6F",X"20",X"50",X"65",X"72",X"65",X"69",X"72",X"61",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 14
		X"20",X"20",X"41",X"6C",X"62",X"65",X"72",X"74",X"6F",X"20",X"4D",X"61",X"69",X"6B",X"75",X"6D",X"61",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 15
		X"20",X"20",X"42",X"72",X"75",X"6E",X"6F",X"20",X"53",X"69",X"6C",X"76",X"61",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 16
		X"20",X"20",X"43",X"61",X"72",X"6C",X"6F",X"73",X"20",X"4B",X"72",X"79",X"6B",X"68",X"74",X"69",X"6E",X"65",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 17
		X"20",X"20",X"43",X"68",X"72",X"69",X"73",X"20",X"48",X"65",X"72",X"62",X"65",X"72",X"74",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 18
		X"20",X"20",X"44",X"2E",X"58",X"61",X"6C",X"69",X"6F",X"72",X"20",X"52",X"69",X"6D",X"72",X"6F",X"6E",X"2D",X"53",X"6F",X"75",X"74",X"74",X"65",X"72",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 19
		X"20",X"20",X"44",X"61",X"76",X"69",X"64",X"20",X"42",X"6F",X"6F",X"63",X"6F",X"63",X"6B",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 20
		X"20",X"20",X"44",X"61",X"76",X"69",X"64",X"20",X"50",X"6F",X"77",X"65",X"6C",X"6C",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 21
		X"20",X"20",X"44",X"61",X"76",X"69",X"64",X"20",X"53",X"61",X"70",X"68",X"69",X"65",X"72",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 22
		X"20",X"20",X"44",X"69",X"6F",X"67",X"6F",X"20",X"50",X"61",X"74",X"72",X"61",X"6F",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 23
		X"20",X"20",X"44",X"69",X"76",X"69",X"6E",X"6F",X"20",X"4C",X"65",X"69",X"74",X"61",X"6F",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 24
		X"20",X"20",X"45",X"64",X"73",X"6F",X"6E",X"20",X"4B",X"61",X"64",X"6F",X"79",X"61",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 25
		X"20",X"20",X"45",X"6D",X"65",X"72",X"73",X"6F",X"6E",X"20",X"43",X"61",X"76",X"61",X"6C",X"6C",X"61",X"72",X"69",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 26
		X"20",X"20",X"47",X"69",X"6C",X"62",X"65",X"72",X"74",X"6F",X"20",X"54",X"61",X"62",X"6F",X"72",X"64",X"61",X"20",X"4A",X"75",X"6E",X"69",X"6F",X"72",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 27
		X"20",X"20",X"48",X"65",X"6E",X"72",X"69",X"71",X"75",X"65",X"20",X"4F",X"6C",X"69",X"66",X"69",X"65",X"72",X"73",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 28
		X"20",X"20",X"48",X"75",X"67",X"6F",X"20",X"47",X"6F",X"6E",X"63",X"61",X"6C",X"76",X"65",X"73",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 29
		X"20",X"20",X"4A",X"6F",X"6E",X"20",X"41",X"72",X"76",X"69",X"64",X"20",X"42",X"6F",X"72",X"72",X"65",X"74",X"7A",X"65",X"6E",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 30
		X"20",X"20",X"4D",X"61",X"6E",X"6F",X"65",X"6C",X"20",X"4C",X"65",X"6D",X"6F",X"73",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 31
		X"20",X"20",X"4D",X"61",X"72",X"69",X"6F",X"20",X"41",X"7A",X"65",X"76",X"65",X"64",X"6F",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 32
		X"20",X"20",X"4D",X"61",X"72",X"63",X"65",X"6C",X"6F",X"20",X"45",X"69",X"72",X"61",X"73",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 33
		X"20",X"20",X"4D",X"61",X"72",X"63",X"65",X"6C",X"6F",X"20",X"46",X"61",X"72",X"69",X"61",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 34
		X"20",X"20",X"4D",X"61",X"72",X"65",X"6B",X"20",X"53",X"7A",X"75",X"6C",X"65",X"6E",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 35
		X"20",X"20",X"4D",X"61",X"72",X"6B",X"20",X"4B",X"6F",X"68",X"6C",X"65",X"72",X"20",X"28",X"4E",X"4D",X"4C",X"33",X"32",X"29",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 36
		X"20",X"20",X"4D",X"61",X"74",X"68",X"65",X"75",X"73",X"20",X"53",X"61",X"6E",X"74",X"6F",X"73",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 37
		X"20",X"20",X"4D",X"61",X"75",X"72",X"6F",X"20",X"50",X"61",X"73",X"73",X"61",X"72",X"69",X"6E",X"68",X"6F",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 38
		X"20",X"20",X"4D",X"61",X"75",X"72",X"69",X"63",X"69",X"6F",X"20",X"41",X"6E",X"64",X"72",X"61",X"64",X"65",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 39
		X"20",X"20",X"4D",X"69",X"6B",X"65",X"20",X"43",X"61",X"64",X"77",X"61",X"6C",X"6C",X"61",X"64",X"65",X"72",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 40
		X"20",X"20",X"50",X"61",X"75",X"6C",X"6F",X"20",X"43",X"61",X"63",X"65",X"6C",X"6C",X"61",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 41
		X"20",X"20",X"50",X"61",X"75",X"6C",X"6F",X"20",X"4D",X"61",X"6C",X"75",X"66",X"20",X"4A",X"72",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 42
		X"20",X"20",X"50",X"65",X"64",X"72",X"6F",X"20",X"4D",X"65",X"64",X"65",X"69",X"72",X"6F",X"73",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 43
		X"20",X"20",X"50",X"61",X"75",X"6C",X"20",X"4C",X"61",X"6E",X"64",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 44
		X"20",X"20",X"50",X"65",X"74",X"65",X"72",X"20",X"46",X"69",X"74",X"63",X"68",X"65",X"74",X"74",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 45
		X"20",X"20",X"50",X"68",X"6F",X"65",X"62",X"75",X"73",X"20",X"44",X"6F",X"6B",X"6F",X"73",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 46
		X"20",X"20",X"52",X"61",X"66",X"61",X"65",X"6C",X"20",X"53",X"69",X"6C",X"76",X"61",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 47
		X"20",X"20",X"52",X"65",X"6E",X"61",X"74",X"6F",X"20",X"47",X"6F",X"6D",X"65",X"73",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 48
		X"20",X"20",X"52",X"6F",X"62",X"65",X"72",X"74",X"20",X"42",X"65",X"72",X"72",X"79",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 49
		X"20",X"20",X"52",X"6F",X"64",X"6F",X"6C",X"66",X"6F",X"20",X"4D",X"61",X"6E",X"6F",X"65",X"6C",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 50
		X"20",X"20",X"52",X"6F",X"6E",X"61",X"6C",X"64",X"6F",X"20",X"50",X"72",X"61",X"64",X"6F",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 51
		X"20",X"20",X"53",X"65",X"76",X"65",X"72",X"69",X"6E",X"6F",X"43",X"76",X"20",X"4A",X"75",X"6E",X"69",X"6F",X"72",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 52
		X"20",X"20",X"54",X"61",X"6D",X"61",X"73",X"20",X"56",X"61",X"6E",X"64",X"6F",X"72",X"66",X"66",X"79",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 53
		X"20",X"20",X"54",X"6F",X"6D",X"20",X"44",X"61",X"6C",X"62",X"79",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 54
		X"20",X"20",X"54",X"6F",X"6E",X"79",X"20",X"55",X"6E",X"64",X"65",X"72",X"77",X"6F",X"6F",X"64",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 55
		X"20",X"20",X"57",X"61",X"6E",X"64",X"65",X"72",X"6C",X"65",X"79",X"20",X"43",X"65",X"73",X"63",X"68",X"69",X"6D",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 56
		X"20",X"20",X"57",X"65",X"72",X"6E",X"65",X"72",X"20",X"4D",X"6F",X"65",X"63",X"6B",X"65",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 57
		X"20",X"20",X"57",X"69",X"6C",X"73",X"6F",X"6E",X"20",X"50",X"69",X"6C",X"6F",X"6E",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 58
		X"20",X"20",X"5A",X"6F",X"6C",X"74",X"61",X"6E",X"20",X"42",X"6F",X"73",X"7A",X"6F",X"72",X"6D",X"65",X"6E",X"79",X"69",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 59
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 60
		X"20",X"20",X"54",X"68",X"61",X"6E",X"6B",X"20",X"79",X"6F",X"75",X"20",X"61",X"6C",X"6C",X"21",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20", -- 61
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20"  -- 62
	);
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
		lines <= x"3f";
	end if;
end process;
end architecture;
