-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80e6",
     9 => x"e4080b0b",
    10 => x"80e6e808",
    11 => x"0b0b80e6",
    12 => x"ec080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"e6ec0c0b",
    16 => x"0b80e6e8",
    17 => x"0c0b0b80",
    18 => x"e6e40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80df9c",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80e6e470",
    57 => x"80f1a027",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c51b192",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80e6",
    65 => x"f40c9f0b",
    66 => x"80e6f80c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"e6f808ff",
    70 => x"0580e6f8",
    71 => x"0c80e6f8",
    72 => x"088025e8",
    73 => x"3880e6f4",
    74 => x"08ff0580",
    75 => x"e6f40c80",
    76 => x"e6f40880",
    77 => x"25d03880",
    78 => x"0b80e6f8",
    79 => x"0c800b80",
    80 => x"e6f40c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80e6f408",
   100 => x"25913882",
   101 => x"c82d80e6",
   102 => x"f408ff05",
   103 => x"80e6f40c",
   104 => x"838a0480",
   105 => x"e6f40880",
   106 => x"e6f80853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80e6f408",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"e6f80881",
   116 => x"0580e6f8",
   117 => x"0c80e6f8",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80e6f8",
   121 => x"0c80e6f4",
   122 => x"08810580",
   123 => x"e6f40c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480e6",
   128 => x"f8088105",
   129 => x"80e6f80c",
   130 => x"80e6f808",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80e6f8",
   134 => x"0c80e6f4",
   135 => x"08810580",
   136 => x"e6f40c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"e6fc0cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"e6fc0c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280e6",
   177 => x"fc088407",
   178 => x"80e6fc0c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b80e3",
   183 => x"b00c8171",
   184 => x"2bff05f6",
   185 => x"880cfdfc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80e6fc",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80e6",
   208 => x"e40c028c",
   209 => x"050d0402",
   210 => x"fc050d81",
   211 => x"808051c0",
   212 => x"115170fb",
   213 => x"38028405",
   214 => x"0d0402fc",
   215 => x"050dec51",
   216 => x"83710c86",
   217 => x"c72d8271",
   218 => x"0c028405",
   219 => x"0d0402fc",
   220 => x"050dec51",
   221 => x"8a710c86",
   222 => x"c72d86c7",
   223 => x"2d86c72d",
   224 => x"86c72d86",
   225 => x"c72d86c7",
   226 => x"2d86c72d",
   227 => x"86c72d86",
   228 => x"c72d86c7",
   229 => x"2d86c72d",
   230 => x"86c72d86",
   231 => x"c72d86c7",
   232 => x"2d86c72d",
   233 => x"86c72d86",
   234 => x"c72d86c7",
   235 => x"2d86c72d",
   236 => x"86c72d86",
   237 => x"c72d86c7",
   238 => x"2d86c72d",
   239 => x"86c72d86",
   240 => x"c72d86c7",
   241 => x"2d86c72d",
   242 => x"86c72d86",
   243 => x"c72d86c7",
   244 => x"2d86c72d",
   245 => x"86c72d86",
   246 => x"c72d86c7",
   247 => x"2d86c72d",
   248 => x"86c72d86",
   249 => x"c72d86c7",
   250 => x"2d86c72d",
   251 => x"86c72d86",
   252 => x"c72d86c7",
   253 => x"2d86c72d",
   254 => x"86c72d86",
   255 => x"c72d86c7",
   256 => x"2d86c72d",
   257 => x"86c72d86",
   258 => x"c72d86c7",
   259 => x"2d86c72d",
   260 => x"86c72d86",
   261 => x"c72d86c7",
   262 => x"2d86c72d",
   263 => x"86c72d86",
   264 => x"c72d86c7",
   265 => x"2d86c72d",
   266 => x"86c72d86",
   267 => x"c72d86c7",
   268 => x"2d86c72d",
   269 => x"86c72d86",
   270 => x"c72d86c7",
   271 => x"2d86c72d",
   272 => x"86c72d86",
   273 => x"c72d86c7",
   274 => x"2d86c72d",
   275 => x"86c72d86",
   276 => x"c72d86c7",
   277 => x"2d86c72d",
   278 => x"86c72d86",
   279 => x"c72d86c7",
   280 => x"2d86c72d",
   281 => x"86c72d86",
   282 => x"c72d86c7",
   283 => x"2d86c72d",
   284 => x"86c72d86",
   285 => x"c72d86c7",
   286 => x"2d86c72d",
   287 => x"86c72d86",
   288 => x"c72d86c7",
   289 => x"2d86c72d",
   290 => x"86c72d86",
   291 => x"c72d86c7",
   292 => x"2d86c72d",
   293 => x"86c72d86",
   294 => x"c72d86c7",
   295 => x"2d86c72d",
   296 => x"86c72d86",
   297 => x"c72d86c7",
   298 => x"2d86c72d",
   299 => x"86c72d86",
   300 => x"c72d86c7",
   301 => x"2d86c72d",
   302 => x"86c72d86",
   303 => x"c72d86c7",
   304 => x"2d86c72d",
   305 => x"86c72d86",
   306 => x"c72d86c7",
   307 => x"2d86c72d",
   308 => x"86c72d86",
   309 => x"c72d86c7",
   310 => x"2d86c72d",
   311 => x"86c72d86",
   312 => x"c72d86c7",
   313 => x"2d86c72d",
   314 => x"86c72d86",
   315 => x"c72d86c7",
   316 => x"2d86c72d",
   317 => x"86c72d86",
   318 => x"c72d86c7",
   319 => x"2d86c72d",
   320 => x"86c72d86",
   321 => x"c72d86c7",
   322 => x"2d86c72d",
   323 => x"86c72d86",
   324 => x"c72d86c7",
   325 => x"2d86c72d",
   326 => x"86c72d86",
   327 => x"c72d86c7",
   328 => x"2d86c72d",
   329 => x"86c72d86",
   330 => x"c72d86c7",
   331 => x"2d86c72d",
   332 => x"86c72d86",
   333 => x"c72d86c7",
   334 => x"2d86c72d",
   335 => x"86c72d86",
   336 => x"c72d86c7",
   337 => x"2d86c72d",
   338 => x"86c72d86",
   339 => x"c72d86c7",
   340 => x"2d86c72d",
   341 => x"86c72d86",
   342 => x"c72d86c7",
   343 => x"2d86c72d",
   344 => x"86c72d86",
   345 => x"c72d86c7",
   346 => x"2d86c72d",
   347 => x"86c72d86",
   348 => x"c72d86c7",
   349 => x"2d86c72d",
   350 => x"86c72d86",
   351 => x"c72d86c7",
   352 => x"2d86c72d",
   353 => x"86c72d86",
   354 => x"c72d86c7",
   355 => x"2d86c72d",
   356 => x"86c72d86",
   357 => x"c72d86c7",
   358 => x"2d86c72d",
   359 => x"86c72d86",
   360 => x"c72d86c7",
   361 => x"2d86c72d",
   362 => x"86c72d86",
   363 => x"c72d86c7",
   364 => x"2d86c72d",
   365 => x"86c72d86",
   366 => x"c72d86c7",
   367 => x"2d86c72d",
   368 => x"86c72d86",
   369 => x"c72d86c7",
   370 => x"2d86c72d",
   371 => x"86c72d86",
   372 => x"c72d86c7",
   373 => x"2d86c72d",
   374 => x"86c72d86",
   375 => x"c72d86c7",
   376 => x"2d86c72d",
   377 => x"86c72d86",
   378 => x"c72d86c7",
   379 => x"2d86c72d",
   380 => x"86c72d86",
   381 => x"c72d86c7",
   382 => x"2d86c72d",
   383 => x"86c72d86",
   384 => x"c72d86c7",
   385 => x"2d86c72d",
   386 => x"86c72d86",
   387 => x"c72d86c7",
   388 => x"2d86c72d",
   389 => x"86c72d86",
   390 => x"c72d86c7",
   391 => x"2d86c72d",
   392 => x"86c72d86",
   393 => x"c72d86c7",
   394 => x"2d86c72d",
   395 => x"86c72d86",
   396 => x"c72d86c7",
   397 => x"2d86c72d",
   398 => x"86c72d86",
   399 => x"c72d86c7",
   400 => x"2d86c72d",
   401 => x"86c72d86",
   402 => x"c72d86c7",
   403 => x"2d86c72d",
   404 => x"86c72d86",
   405 => x"c72d86c7",
   406 => x"2d86c72d",
   407 => x"86c72d86",
   408 => x"c72d86c7",
   409 => x"2d86c72d",
   410 => x"86c72d86",
   411 => x"c72d86c7",
   412 => x"2d86c72d",
   413 => x"86c72d86",
   414 => x"c72d86c7",
   415 => x"2d86c72d",
   416 => x"86c72d86",
   417 => x"c72d86c7",
   418 => x"2d86c72d",
   419 => x"86c72d86",
   420 => x"c72d86c7",
   421 => x"2d86c72d",
   422 => x"86c72d86",
   423 => x"c72d86c7",
   424 => x"2d86c72d",
   425 => x"86c72d86",
   426 => x"c72d86c7",
   427 => x"2d86c72d",
   428 => x"86c72d86",
   429 => x"c72d86c7",
   430 => x"2d86c72d",
   431 => x"86c72d86",
   432 => x"c72d86c7",
   433 => x"2d86c72d",
   434 => x"86c72d86",
   435 => x"c72d86c7",
   436 => x"2d86c72d",
   437 => x"86c72d86",
   438 => x"c72d86c7",
   439 => x"2d86c72d",
   440 => x"86c72d86",
   441 => x"c72d86c7",
   442 => x"2d86c72d",
   443 => x"86c72d86",
   444 => x"c72d86c7",
   445 => x"2d86c72d",
   446 => x"86c72d86",
   447 => x"c72d86c7",
   448 => x"2d86c72d",
   449 => x"86c72d86",
   450 => x"c72d86c7",
   451 => x"2d86c72d",
   452 => x"86c72d86",
   453 => x"c72d86c7",
   454 => x"2d86c72d",
   455 => x"86c72d86",
   456 => x"c72d86c7",
   457 => x"2d86c72d",
   458 => x"86c72d86",
   459 => x"c72d86c7",
   460 => x"2d86c72d",
   461 => x"86c72d86",
   462 => x"c72d86c7",
   463 => x"2d86c72d",
   464 => x"86c72d86",
   465 => x"c72d86c7",
   466 => x"2d86c72d",
   467 => x"86c72d86",
   468 => x"c72d86c7",
   469 => x"2d86c72d",
   470 => x"86c72d86",
   471 => x"c72d86c7",
   472 => x"2d86c72d",
   473 => x"86c72d86",
   474 => x"c72d86c7",
   475 => x"2d86c72d",
   476 => x"86c72d86",
   477 => x"c72d86c7",
   478 => x"2d86c72d",
   479 => x"86c72d86",
   480 => x"c72d86c7",
   481 => x"2d86c72d",
   482 => x"86c72d86",
   483 => x"c72d86c7",
   484 => x"2d86c72d",
   485 => x"86c72d86",
   486 => x"c72d86c7",
   487 => x"2d86c72d",
   488 => x"86c72d86",
   489 => x"c72d86c7",
   490 => x"2d86c72d",
   491 => x"86c72d86",
   492 => x"c72d86c7",
   493 => x"2d86c72d",
   494 => x"86c72d86",
   495 => x"c72d86c7",
   496 => x"2d86c72d",
   497 => x"86c72d86",
   498 => x"c72d86c7",
   499 => x"2d86c72d",
   500 => x"86c72d86",
   501 => x"c72d86c7",
   502 => x"2d86c72d",
   503 => x"86c72d86",
   504 => x"c72d86c7",
   505 => x"2d86c72d",
   506 => x"86c72d86",
   507 => x"c72d86c7",
   508 => x"2d86c72d",
   509 => x"86c72d86",
   510 => x"c72d86c7",
   511 => x"2d86c72d",
   512 => x"86c72d86",
   513 => x"c72d86c7",
   514 => x"2d86c72d",
   515 => x"86c72d86",
   516 => x"c72d86c7",
   517 => x"2d86c72d",
   518 => x"86c72d86",
   519 => x"c72d86c7",
   520 => x"2d86c72d",
   521 => x"86c72d86",
   522 => x"c72d86c7",
   523 => x"2d86c72d",
   524 => x"86c72d86",
   525 => x"c72d86c7",
   526 => x"2d86c72d",
   527 => x"86c72d86",
   528 => x"c72d86c7",
   529 => x"2d86c72d",
   530 => x"86c72d86",
   531 => x"c72d86c7",
   532 => x"2d86c72d",
   533 => x"86c72d86",
   534 => x"c72d86c7",
   535 => x"2d86c72d",
   536 => x"86c72d86",
   537 => x"c72d86c7",
   538 => x"2d86c72d",
   539 => x"86c72d86",
   540 => x"c72d86c7",
   541 => x"2d86c72d",
   542 => x"86c72d86",
   543 => x"c72d86c7",
   544 => x"2d86c72d",
   545 => x"86c72d86",
   546 => x"c72d86c7",
   547 => x"2d86c72d",
   548 => x"86c72d86",
   549 => x"c72d86c7",
   550 => x"2d86c72d",
   551 => x"86c72d86",
   552 => x"c72d86c7",
   553 => x"2d86c72d",
   554 => x"86c72d86",
   555 => x"c72d86c7",
   556 => x"2d86c72d",
   557 => x"86c72d86",
   558 => x"c72d86c7",
   559 => x"2d86c72d",
   560 => x"86c72d86",
   561 => x"c72d86c7",
   562 => x"2d86c72d",
   563 => x"86c72d86",
   564 => x"c72d86c7",
   565 => x"2d86c72d",
   566 => x"86c72d86",
   567 => x"c72d86c7",
   568 => x"2d86c72d",
   569 => x"86c72d86",
   570 => x"c72d86c7",
   571 => x"2d86c72d",
   572 => x"86c72d86",
   573 => x"c72d86c7",
   574 => x"2d86c72d",
   575 => x"86c72d86",
   576 => x"c72d86c7",
   577 => x"2d86c72d",
   578 => x"86c72d86",
   579 => x"c72d86c7",
   580 => x"2d86c72d",
   581 => x"86c72d86",
   582 => x"c72d86c7",
   583 => x"2d86c72d",
   584 => x"86c72d86",
   585 => x"c72d86c7",
   586 => x"2d86c72d",
   587 => x"86c72d86",
   588 => x"c72d86c7",
   589 => x"2d86c72d",
   590 => x"86c72d86",
   591 => x"c72d86c7",
   592 => x"2d86c72d",
   593 => x"86c72d86",
   594 => x"c72d86c7",
   595 => x"2d86c72d",
   596 => x"86c72d86",
   597 => x"c72d86c7",
   598 => x"2d86c72d",
   599 => x"86c72d86",
   600 => x"c72d86c7",
   601 => x"2d86c72d",
   602 => x"86c72d86",
   603 => x"c72d86c7",
   604 => x"2d86c72d",
   605 => x"86c72d86",
   606 => x"c72d86c7",
   607 => x"2d86c72d",
   608 => x"86c72d86",
   609 => x"c72d86c7",
   610 => x"2d86c72d",
   611 => x"86c72d86",
   612 => x"c72d86c7",
   613 => x"2d86c72d",
   614 => x"86c72d86",
   615 => x"c72d86c7",
   616 => x"2d86c72d",
   617 => x"86c72d86",
   618 => x"c72d86c7",
   619 => x"2d86c72d",
   620 => x"86c72d86",
   621 => x"c72d86c7",
   622 => x"2d86c72d",
   623 => x"86c72d86",
   624 => x"c72d86c7",
   625 => x"2d86c72d",
   626 => x"86c72d86",
   627 => x"c72d86c7",
   628 => x"2d86c72d",
   629 => x"86c72d86",
   630 => x"c72d86c7",
   631 => x"2d86c72d",
   632 => x"86c72d86",
   633 => x"c72d86c7",
   634 => x"2d86c72d",
   635 => x"86c72d86",
   636 => x"c72d86c7",
   637 => x"2d86c72d",
   638 => x"86c72d86",
   639 => x"c72d86c7",
   640 => x"2d86c72d",
   641 => x"86c72d86",
   642 => x"c72d86c7",
   643 => x"2d86c72d",
   644 => x"86c72d86",
   645 => x"c72d86c7",
   646 => x"2d86c72d",
   647 => x"86c72d86",
   648 => x"c72d86c7",
   649 => x"2d86c72d",
   650 => x"86c72d86",
   651 => x"c72d86c7",
   652 => x"2d86c72d",
   653 => x"86c72d82",
   654 => x"710c0284",
   655 => x"050d0402",
   656 => x"fc050dec",
   657 => x"5192710c",
   658 => x"86c72d86",
   659 => x"c72d86c7",
   660 => x"2d86c72d",
   661 => x"86c72d86",
   662 => x"c72d86c7",
   663 => x"2d86c72d",
   664 => x"86c72d86",
   665 => x"c72d86c7",
   666 => x"2d86c72d",
   667 => x"86c72d86",
   668 => x"c72d86c7",
   669 => x"2d86c72d",
   670 => x"86c72d86",
   671 => x"c72d86c7",
   672 => x"2d86c72d",
   673 => x"86c72d86",
   674 => x"c72d86c7",
   675 => x"2d86c72d",
   676 => x"86c72d86",
   677 => x"c72d86c7",
   678 => x"2d86c72d",
   679 => x"86c72d86",
   680 => x"c72d86c7",
   681 => x"2d86c72d",
   682 => x"86c72d86",
   683 => x"c72d86c7",
   684 => x"2d86c72d",
   685 => x"86c72d86",
   686 => x"c72d86c7",
   687 => x"2d86c72d",
   688 => x"86c72d86",
   689 => x"c72d86c7",
   690 => x"2d86c72d",
   691 => x"86c72d86",
   692 => x"c72d86c7",
   693 => x"2d86c72d",
   694 => x"86c72d86",
   695 => x"c72d86c7",
   696 => x"2d86c72d",
   697 => x"86c72d86",
   698 => x"c72d86c7",
   699 => x"2d86c72d",
   700 => x"86c72d86",
   701 => x"c72d86c7",
   702 => x"2d86c72d",
   703 => x"86c72d86",
   704 => x"c72d86c7",
   705 => x"2d86c72d",
   706 => x"86c72d86",
   707 => x"c72d86c7",
   708 => x"2d86c72d",
   709 => x"86c72d86",
   710 => x"c72d86c7",
   711 => x"2d86c72d",
   712 => x"86c72d86",
   713 => x"c72d86c7",
   714 => x"2d86c72d",
   715 => x"86c72d86",
   716 => x"c72d86c7",
   717 => x"2d86c72d",
   718 => x"86c72d86",
   719 => x"c72d86c7",
   720 => x"2d86c72d",
   721 => x"86c72d86",
   722 => x"c72d86c7",
   723 => x"2d86c72d",
   724 => x"86c72d86",
   725 => x"c72d86c7",
   726 => x"2d86c72d",
   727 => x"86c72d86",
   728 => x"c72d86c7",
   729 => x"2d86c72d",
   730 => x"86c72d86",
   731 => x"c72d86c7",
   732 => x"2d86c72d",
   733 => x"86c72d86",
   734 => x"c72d86c7",
   735 => x"2d86c72d",
   736 => x"86c72d86",
   737 => x"c72d86c7",
   738 => x"2d86c72d",
   739 => x"86c72d86",
   740 => x"c72d86c7",
   741 => x"2d86c72d",
   742 => x"86c72d86",
   743 => x"c72d86c7",
   744 => x"2d86c72d",
   745 => x"86c72d86",
   746 => x"c72d86c7",
   747 => x"2d86c72d",
   748 => x"86c72d86",
   749 => x"c72d86c7",
   750 => x"2d86c72d",
   751 => x"86c72d86",
   752 => x"c72d86c7",
   753 => x"2d86c72d",
   754 => x"86c72d86",
   755 => x"c72d86c7",
   756 => x"2d86c72d",
   757 => x"86c72d86",
   758 => x"c72d86c7",
   759 => x"2d86c72d",
   760 => x"86c72d86",
   761 => x"c72d86c7",
   762 => x"2d86c72d",
   763 => x"86c72d86",
   764 => x"c72d86c7",
   765 => x"2d86c72d",
   766 => x"86c72d86",
   767 => x"c72d86c7",
   768 => x"2d86c72d",
   769 => x"86c72d86",
   770 => x"c72d86c7",
   771 => x"2d86c72d",
   772 => x"86c72d86",
   773 => x"c72d86c7",
   774 => x"2d86c72d",
   775 => x"86c72d86",
   776 => x"c72d86c7",
   777 => x"2d86c72d",
   778 => x"86c72d86",
   779 => x"c72d86c7",
   780 => x"2d86c72d",
   781 => x"86c72d86",
   782 => x"c72d86c7",
   783 => x"2d86c72d",
   784 => x"86c72d86",
   785 => x"c72d86c7",
   786 => x"2d86c72d",
   787 => x"86c72d86",
   788 => x"c72d86c7",
   789 => x"2d86c72d",
   790 => x"86c72d86",
   791 => x"c72d86c7",
   792 => x"2d86c72d",
   793 => x"86c72d86",
   794 => x"c72d86c7",
   795 => x"2d86c72d",
   796 => x"86c72d86",
   797 => x"c72d86c7",
   798 => x"2d86c72d",
   799 => x"86c72d86",
   800 => x"c72d86c7",
   801 => x"2d86c72d",
   802 => x"86c72d86",
   803 => x"c72d86c7",
   804 => x"2d86c72d",
   805 => x"86c72d86",
   806 => x"c72d86c7",
   807 => x"2d86c72d",
   808 => x"86c72d86",
   809 => x"c72d86c7",
   810 => x"2d86c72d",
   811 => x"86c72d86",
   812 => x"c72d86c7",
   813 => x"2d86c72d",
   814 => x"86c72d86",
   815 => x"c72d86c7",
   816 => x"2d86c72d",
   817 => x"86c72d86",
   818 => x"c72d86c7",
   819 => x"2d86c72d",
   820 => x"86c72d86",
   821 => x"c72d86c7",
   822 => x"2d86c72d",
   823 => x"86c72d86",
   824 => x"c72d86c7",
   825 => x"2d86c72d",
   826 => x"86c72d86",
   827 => x"c72d86c7",
   828 => x"2d86c72d",
   829 => x"86c72d86",
   830 => x"c72d86c7",
   831 => x"2d86c72d",
   832 => x"86c72d86",
   833 => x"c72d86c7",
   834 => x"2d86c72d",
   835 => x"86c72d86",
   836 => x"c72d86c7",
   837 => x"2d86c72d",
   838 => x"86c72d86",
   839 => x"c72d86c7",
   840 => x"2d86c72d",
   841 => x"86c72d86",
   842 => x"c72d86c7",
   843 => x"2d86c72d",
   844 => x"86c72d86",
   845 => x"c72d86c7",
   846 => x"2d86c72d",
   847 => x"86c72d86",
   848 => x"c72d86c7",
   849 => x"2d86c72d",
   850 => x"86c72d86",
   851 => x"c72d86c7",
   852 => x"2d86c72d",
   853 => x"86c72d86",
   854 => x"c72d86c7",
   855 => x"2d86c72d",
   856 => x"86c72d86",
   857 => x"c72d86c7",
   858 => x"2d86c72d",
   859 => x"86c72d86",
   860 => x"c72d86c7",
   861 => x"2d86c72d",
   862 => x"86c72d86",
   863 => x"c72d86c7",
   864 => x"2d86c72d",
   865 => x"86c72d86",
   866 => x"c72d86c7",
   867 => x"2d86c72d",
   868 => x"86c72d86",
   869 => x"c72d86c7",
   870 => x"2d86c72d",
   871 => x"86c72d86",
   872 => x"c72d86c7",
   873 => x"2d86c72d",
   874 => x"86c72d86",
   875 => x"c72d86c7",
   876 => x"2d86c72d",
   877 => x"86c72d86",
   878 => x"c72d86c7",
   879 => x"2d86c72d",
   880 => x"86c72d86",
   881 => x"c72d86c7",
   882 => x"2d86c72d",
   883 => x"86c72d86",
   884 => x"c72d86c7",
   885 => x"2d86c72d",
   886 => x"86c72d86",
   887 => x"c72d86c7",
   888 => x"2d86c72d",
   889 => x"86c72d86",
   890 => x"c72d86c7",
   891 => x"2d86c72d",
   892 => x"86c72d86",
   893 => x"c72d86c7",
   894 => x"2d86c72d",
   895 => x"86c72d86",
   896 => x"c72d86c7",
   897 => x"2d86c72d",
   898 => x"86c72d86",
   899 => x"c72d86c7",
   900 => x"2d86c72d",
   901 => x"86c72d86",
   902 => x"c72d86c7",
   903 => x"2d86c72d",
   904 => x"86c72d86",
   905 => x"c72d86c7",
   906 => x"2d86c72d",
   907 => x"86c72d86",
   908 => x"c72d86c7",
   909 => x"2d86c72d",
   910 => x"86c72d86",
   911 => x"c72d86c7",
   912 => x"2d86c72d",
   913 => x"86c72d86",
   914 => x"c72d86c7",
   915 => x"2d86c72d",
   916 => x"86c72d86",
   917 => x"c72d86c7",
   918 => x"2d86c72d",
   919 => x"86c72d86",
   920 => x"c72d86c7",
   921 => x"2d86c72d",
   922 => x"86c72d86",
   923 => x"c72d86c7",
   924 => x"2d86c72d",
   925 => x"86c72d86",
   926 => x"c72d86c7",
   927 => x"2d86c72d",
   928 => x"86c72d86",
   929 => x"c72d86c7",
   930 => x"2d86c72d",
   931 => x"86c72d86",
   932 => x"c72d86c7",
   933 => x"2d86c72d",
   934 => x"86c72d86",
   935 => x"c72d86c7",
   936 => x"2d86c72d",
   937 => x"86c72d86",
   938 => x"c72d86c7",
   939 => x"2d86c72d",
   940 => x"86c72d86",
   941 => x"c72d86c7",
   942 => x"2d86c72d",
   943 => x"86c72d86",
   944 => x"c72d86c7",
   945 => x"2d86c72d",
   946 => x"86c72d86",
   947 => x"c72d86c7",
   948 => x"2d86c72d",
   949 => x"86c72d86",
   950 => x"c72d86c7",
   951 => x"2d86c72d",
   952 => x"86c72d86",
   953 => x"c72d86c7",
   954 => x"2d86c72d",
   955 => x"86c72d86",
   956 => x"c72d86c7",
   957 => x"2d86c72d",
   958 => x"86c72d86",
   959 => x"c72d86c7",
   960 => x"2d86c72d",
   961 => x"86c72d86",
   962 => x"c72d86c7",
   963 => x"2d86c72d",
   964 => x"86c72d86",
   965 => x"c72d86c7",
   966 => x"2d86c72d",
   967 => x"86c72d86",
   968 => x"c72d86c7",
   969 => x"2d86c72d",
   970 => x"86c72d86",
   971 => x"c72d86c7",
   972 => x"2d86c72d",
   973 => x"86c72d86",
   974 => x"c72d86c7",
   975 => x"2d86c72d",
   976 => x"86c72d86",
   977 => x"c72d86c7",
   978 => x"2d86c72d",
   979 => x"86c72d86",
   980 => x"c72d86c7",
   981 => x"2d86c72d",
   982 => x"86c72d86",
   983 => x"c72d86c7",
   984 => x"2d86c72d",
   985 => x"86c72d86",
   986 => x"c72d86c7",
   987 => x"2d86c72d",
   988 => x"86c72d86",
   989 => x"c72d86c7",
   990 => x"2d86c72d",
   991 => x"86c72d86",
   992 => x"c72d86c7",
   993 => x"2d86c72d",
   994 => x"86c72d86",
   995 => x"c72d86c7",
   996 => x"2d86c72d",
   997 => x"86c72d86",
   998 => x"c72d86c7",
   999 => x"2d86c72d",
  1000 => x"86c72d86",
  1001 => x"c72d86c7",
  1002 => x"2d86c72d",
  1003 => x"86c72d86",
  1004 => x"c72d86c7",
  1005 => x"2d86c72d",
  1006 => x"86c72d86",
  1007 => x"c72d86c7",
  1008 => x"2d86c72d",
  1009 => x"86c72d86",
  1010 => x"c72d86c7",
  1011 => x"2d86c72d",
  1012 => x"86c72d86",
  1013 => x"c72d86c7",
  1014 => x"2d86c72d",
  1015 => x"86c72d86",
  1016 => x"c72d86c7",
  1017 => x"2d86c72d",
  1018 => x"86c72d86",
  1019 => x"c72d86c7",
  1020 => x"2d86c72d",
  1021 => x"86c72d86",
  1022 => x"c72d86c7",
  1023 => x"2d86c72d",
  1024 => x"86c72d86",
  1025 => x"c72d86c7",
  1026 => x"2d86c72d",
  1027 => x"86c72d86",
  1028 => x"c72d86c7",
  1029 => x"2d86c72d",
  1030 => x"86c72d86",
  1031 => x"c72d86c7",
  1032 => x"2d86c72d",
  1033 => x"86c72d86",
  1034 => x"c72d86c7",
  1035 => x"2d86c72d",
  1036 => x"86c72d86",
  1037 => x"c72d86c7",
  1038 => x"2d86c72d",
  1039 => x"86c72d86",
  1040 => x"c72d86c7",
  1041 => x"2d86c72d",
  1042 => x"86c72d86",
  1043 => x"c72d86c7",
  1044 => x"2d86c72d",
  1045 => x"86c72d86",
  1046 => x"c72d86c7",
  1047 => x"2d86c72d",
  1048 => x"86c72d86",
  1049 => x"c72d86c7",
  1050 => x"2d86c72d",
  1051 => x"86c72d86",
  1052 => x"c72d86c7",
  1053 => x"2d86c72d",
  1054 => x"86c72d86",
  1055 => x"c72d86c7",
  1056 => x"2d86c72d",
  1057 => x"86c72d86",
  1058 => x"c72d86c7",
  1059 => x"2d86c72d",
  1060 => x"86c72d86",
  1061 => x"c72d86c7",
  1062 => x"2d86c72d",
  1063 => x"86c72d86",
  1064 => x"c72d86c7",
  1065 => x"2d86c72d",
  1066 => x"86c72d86",
  1067 => x"c72d86c7",
  1068 => x"2d86c72d",
  1069 => x"86c72d86",
  1070 => x"c72d86c7",
  1071 => x"2d86c72d",
  1072 => x"86c72d86",
  1073 => x"c72d86c7",
  1074 => x"2d86c72d",
  1075 => x"86c72d86",
  1076 => x"c72d86c7",
  1077 => x"2d86c72d",
  1078 => x"86c72d86",
  1079 => x"c72d86c7",
  1080 => x"2d86c72d",
  1081 => x"86c72d86",
  1082 => x"c72d86c7",
  1083 => x"2d86c72d",
  1084 => x"86c72d86",
  1085 => x"c72d86c7",
  1086 => x"2d86c72d",
  1087 => x"86c72d86",
  1088 => x"c72d86c7",
  1089 => x"2d86c72d",
  1090 => x"82710c02",
  1091 => x"84050d04",
  1092 => x"a00bec0c",
  1093 => x"86c72d86",
  1094 => x"c72d86c7",
  1095 => x"2d86c72d",
  1096 => x"86c72d86",
  1097 => x"c72d86c7",
  1098 => x"2d86c72d",
  1099 => x"86c72d86",
  1100 => x"c72d86c7",
  1101 => x"2d86c72d",
  1102 => x"86c72d86",
  1103 => x"c72d86c7",
  1104 => x"2d86c72d",
  1105 => x"86c72d86",
  1106 => x"c72d86c7",
  1107 => x"2d86c72d",
  1108 => x"86c72d86",
  1109 => x"c72d86c7",
  1110 => x"2d86c72d",
  1111 => x"86c72d86",
  1112 => x"c72d86c7",
  1113 => x"2d86c72d",
  1114 => x"86c72d86",
  1115 => x"c72d86c7",
  1116 => x"2d86c72d",
  1117 => x"86c72d86",
  1118 => x"c72d86c7",
  1119 => x"2d86c72d",
  1120 => x"86c72d86",
  1121 => x"c72d86c7",
  1122 => x"2d86c72d",
  1123 => x"86c72d86",
  1124 => x"c72d86c7",
  1125 => x"2d86c72d",
  1126 => x"86c72d86",
  1127 => x"c72d86c7",
  1128 => x"2d86c72d",
  1129 => x"86c72d86",
  1130 => x"c72d86c7",
  1131 => x"2d86c72d",
  1132 => x"86c72d86",
  1133 => x"c72d86c7",
  1134 => x"2d86c72d",
  1135 => x"86c72d86",
  1136 => x"c72d86c7",
  1137 => x"2d86c72d",
  1138 => x"86c72d86",
  1139 => x"c72d86c7",
  1140 => x"2d86c72d",
  1141 => x"86c72d86",
  1142 => x"c72d86c7",
  1143 => x"2d86c72d",
  1144 => x"86c72d86",
  1145 => x"c72d86c7",
  1146 => x"2d86c72d",
  1147 => x"86c72d86",
  1148 => x"c72d86c7",
  1149 => x"2d86c72d",
  1150 => x"86c72d86",
  1151 => x"c72d86c7",
  1152 => x"2d86c72d",
  1153 => x"86c72d86",
  1154 => x"c72d86c7",
  1155 => x"2d86c72d",
  1156 => x"86c72d86",
  1157 => x"c72d86c7",
  1158 => x"2d86c72d",
  1159 => x"86c72d86",
  1160 => x"c72d86c7",
  1161 => x"2d86c72d",
  1162 => x"86c72d86",
  1163 => x"c72d86c7",
  1164 => x"2d86c72d",
  1165 => x"86c72d86",
  1166 => x"c72d86c7",
  1167 => x"2d86c72d",
  1168 => x"86c72d86",
  1169 => x"c72d86c7",
  1170 => x"2d86c72d",
  1171 => x"86c72d86",
  1172 => x"c72d86c7",
  1173 => x"2d86c72d",
  1174 => x"86c72d86",
  1175 => x"c72d86c7",
  1176 => x"2d86c72d",
  1177 => x"86c72d86",
  1178 => x"c72d86c7",
  1179 => x"2d86c72d",
  1180 => x"86c72d86",
  1181 => x"c72d86c7",
  1182 => x"2d86c72d",
  1183 => x"86c72d86",
  1184 => x"c72d86c7",
  1185 => x"2d86c72d",
  1186 => x"86c72d86",
  1187 => x"c72d86c7",
  1188 => x"2d86c72d",
  1189 => x"86c72d86",
  1190 => x"c72d86c7",
  1191 => x"2d86c72d",
  1192 => x"86c72d86",
  1193 => x"c72d86c7",
  1194 => x"2d86c72d",
  1195 => x"86c72d86",
  1196 => x"c72d86c7",
  1197 => x"2d86c72d",
  1198 => x"86c72d86",
  1199 => x"c72d86c7",
  1200 => x"2d86c72d",
  1201 => x"86c72d86",
  1202 => x"c72d86c7",
  1203 => x"2d86c72d",
  1204 => x"86c72d86",
  1205 => x"c72d86c7",
  1206 => x"2d86c72d",
  1207 => x"86c72d86",
  1208 => x"c72d86c7",
  1209 => x"2d86c72d",
  1210 => x"86c72d86",
  1211 => x"c72d86c7",
  1212 => x"2d86c72d",
  1213 => x"86c72d86",
  1214 => x"c72d86c7",
  1215 => x"2d86c72d",
  1216 => x"86c72d86",
  1217 => x"c72d86c7",
  1218 => x"2d86c72d",
  1219 => x"86c72d86",
  1220 => x"c72d86c7",
  1221 => x"2d86c72d",
  1222 => x"86c72d86",
  1223 => x"c72d86c7",
  1224 => x"2d86c72d",
  1225 => x"86c72d86",
  1226 => x"c72d86c7",
  1227 => x"2d86c72d",
  1228 => x"86c72d86",
  1229 => x"c72d86c7",
  1230 => x"2d86c72d",
  1231 => x"86c72d86",
  1232 => x"c72d86c7",
  1233 => x"2d86c72d",
  1234 => x"86c72d86",
  1235 => x"c72d86c7",
  1236 => x"2d86c72d",
  1237 => x"86c72d86",
  1238 => x"c72d86c7",
  1239 => x"2d86c72d",
  1240 => x"86c72d86",
  1241 => x"c72d86c7",
  1242 => x"2d86c72d",
  1243 => x"86c72d86",
  1244 => x"c72d86c7",
  1245 => x"2d86c72d",
  1246 => x"86c72d86",
  1247 => x"c72d86c7",
  1248 => x"2d86c72d",
  1249 => x"86c72d86",
  1250 => x"c72d86c7",
  1251 => x"2d86c72d",
  1252 => x"86c72d86",
  1253 => x"c72d86c7",
  1254 => x"2d86c72d",
  1255 => x"86c72d86",
  1256 => x"c72d86c7",
  1257 => x"2d86c72d",
  1258 => x"86c72d86",
  1259 => x"c72d86c7",
  1260 => x"2d86c72d",
  1261 => x"86c72d86",
  1262 => x"c72d86c7",
  1263 => x"2d86c72d",
  1264 => x"86c72d86",
  1265 => x"c72d86c7",
  1266 => x"2d86c72d",
  1267 => x"86c72d86",
  1268 => x"c72d86c7",
  1269 => x"2d86c72d",
  1270 => x"86c72d86",
  1271 => x"c72d86c7",
  1272 => x"2d86c72d",
  1273 => x"86c72d86",
  1274 => x"c72d86c7",
  1275 => x"2d86c72d",
  1276 => x"86c72d86",
  1277 => x"c72d86c7",
  1278 => x"2d86c72d",
  1279 => x"86c72d86",
  1280 => x"c72d86c7",
  1281 => x"2d86c72d",
  1282 => x"86c72d86",
  1283 => x"c72d86c7",
  1284 => x"2d86c72d",
  1285 => x"86c72d86",
  1286 => x"c72d86c7",
  1287 => x"2d86c72d",
  1288 => x"86c72d86",
  1289 => x"c72d86c7",
  1290 => x"2d86c72d",
  1291 => x"86c72d86",
  1292 => x"c72d86c7",
  1293 => x"2d86c72d",
  1294 => x"86c72d86",
  1295 => x"c72d86c7",
  1296 => x"2d86c72d",
  1297 => x"86c72d86",
  1298 => x"c72d86c7",
  1299 => x"2d86c72d",
  1300 => x"86c72d86",
  1301 => x"c72d86c7",
  1302 => x"2d86c72d",
  1303 => x"86c72d86",
  1304 => x"c72d86c7",
  1305 => x"2d86c72d",
  1306 => x"86c72d86",
  1307 => x"c72d86c7",
  1308 => x"2d86c72d",
  1309 => x"86c72d86",
  1310 => x"c72d86c7",
  1311 => x"2d86c72d",
  1312 => x"86c72d86",
  1313 => x"c72d86c7",
  1314 => x"2d86c72d",
  1315 => x"86c72d86",
  1316 => x"c72d86c7",
  1317 => x"2d86c72d",
  1318 => x"86c72d86",
  1319 => x"c72d86c7",
  1320 => x"2d86c72d",
  1321 => x"86c72d86",
  1322 => x"c72d86c7",
  1323 => x"2d86c72d",
  1324 => x"86c72d86",
  1325 => x"c72d86c7",
  1326 => x"2d86c72d",
  1327 => x"86c72d86",
  1328 => x"c72d86c7",
  1329 => x"2d86c72d",
  1330 => x"86c72d86",
  1331 => x"c72d86c7",
  1332 => x"2d86c72d",
  1333 => x"86c72d86",
  1334 => x"c72d86c7",
  1335 => x"2d86c72d",
  1336 => x"86c72d86",
  1337 => x"c72d86c7",
  1338 => x"2d86c72d",
  1339 => x"86c72d86",
  1340 => x"c72d86c7",
  1341 => x"2d86c72d",
  1342 => x"86c72d86",
  1343 => x"c72d86c7",
  1344 => x"2d86c72d",
  1345 => x"86c72d86",
  1346 => x"c72d86c7",
  1347 => x"2d86c72d",
  1348 => x"86c72d86",
  1349 => x"c72d86c7",
  1350 => x"2d86c72d",
  1351 => x"86c72d86",
  1352 => x"c72d86c7",
  1353 => x"2d86c72d",
  1354 => x"86c72d86",
  1355 => x"c72d86c7",
  1356 => x"2d86c72d",
  1357 => x"86c72d86",
  1358 => x"c72d86c7",
  1359 => x"2d86c72d",
  1360 => x"86c72d86",
  1361 => x"c72d86c7",
  1362 => x"2d86c72d",
  1363 => x"86c72d86",
  1364 => x"c72d86c7",
  1365 => x"2d86c72d",
  1366 => x"86c72d86",
  1367 => x"c72d86c7",
  1368 => x"2d86c72d",
  1369 => x"86c72d86",
  1370 => x"c72d86c7",
  1371 => x"2d86c72d",
  1372 => x"86c72d86",
  1373 => x"c72d86c7",
  1374 => x"2d86c72d",
  1375 => x"86c72d86",
  1376 => x"c72d86c7",
  1377 => x"2d86c72d",
  1378 => x"86c72d86",
  1379 => x"c72d86c7",
  1380 => x"2d86c72d",
  1381 => x"86c72d86",
  1382 => x"c72d86c7",
  1383 => x"2d86c72d",
  1384 => x"86c72d86",
  1385 => x"c72d86c7",
  1386 => x"2d86c72d",
  1387 => x"86c72d86",
  1388 => x"c72d86c7",
  1389 => x"2d86c72d",
  1390 => x"86c72d86",
  1391 => x"c72d86c7",
  1392 => x"2d86c72d",
  1393 => x"86c72d86",
  1394 => x"c72d86c7",
  1395 => x"2d86c72d",
  1396 => x"86c72d86",
  1397 => x"c72d86c7",
  1398 => x"2d86c72d",
  1399 => x"86c72d86",
  1400 => x"c72d86c7",
  1401 => x"2d86c72d",
  1402 => x"86c72d86",
  1403 => x"c72d86c7",
  1404 => x"2d86c72d",
  1405 => x"86c72d86",
  1406 => x"c72d86c7",
  1407 => x"2d86c72d",
  1408 => x"86c72d86",
  1409 => x"c72d86c7",
  1410 => x"2d86c72d",
  1411 => x"86c72d86",
  1412 => x"c72d86c7",
  1413 => x"2d86c72d",
  1414 => x"86c72d86",
  1415 => x"c72d86c7",
  1416 => x"2d86c72d",
  1417 => x"86c72d86",
  1418 => x"c72d86c7",
  1419 => x"2d86c72d",
  1420 => x"86c72d86",
  1421 => x"c72d86c7",
  1422 => x"2d86c72d",
  1423 => x"86c72d86",
  1424 => x"c72d86c7",
  1425 => x"2d86c72d",
  1426 => x"86c72d86",
  1427 => x"c72d86c7",
  1428 => x"2d86c72d",
  1429 => x"86c72d86",
  1430 => x"c72d86c7",
  1431 => x"2d86c72d",
  1432 => x"86c72d86",
  1433 => x"c72d86c7",
  1434 => x"2d86c72d",
  1435 => x"86c72d86",
  1436 => x"c72d86c7",
  1437 => x"2d86c72d",
  1438 => x"86c72d86",
  1439 => x"c72d86c7",
  1440 => x"2d86c72d",
  1441 => x"86c72d86",
  1442 => x"c72d86c7",
  1443 => x"2d86c72d",
  1444 => x"86c72d86",
  1445 => x"c72d86c7",
  1446 => x"2d86c72d",
  1447 => x"86c72d86",
  1448 => x"c72d86c7",
  1449 => x"2d86c72d",
  1450 => x"86c72d86",
  1451 => x"c72d86c7",
  1452 => x"2d86c72d",
  1453 => x"86c72d86",
  1454 => x"c72d86c7",
  1455 => x"2d86c72d",
  1456 => x"86c72d86",
  1457 => x"c72d86c7",
  1458 => x"2d86c72d",
  1459 => x"86c72d86",
  1460 => x"c72d86c7",
  1461 => x"2d86c72d",
  1462 => x"86c72d86",
  1463 => x"c72d86c7",
  1464 => x"2d86c72d",
  1465 => x"86c72d86",
  1466 => x"c72d86c7",
  1467 => x"2d86c72d",
  1468 => x"86c72d86",
  1469 => x"c72d86c7",
  1470 => x"2d86c72d",
  1471 => x"86c72d86",
  1472 => x"c72d86c7",
  1473 => x"2d86c72d",
  1474 => x"86c72d86",
  1475 => x"c72d86c7",
  1476 => x"2d86c72d",
  1477 => x"86c72d86",
  1478 => x"c72d86c7",
  1479 => x"2d86c72d",
  1480 => x"86c72d86",
  1481 => x"c72d86c7",
  1482 => x"2d86c72d",
  1483 => x"86c72d86",
  1484 => x"c72d86c7",
  1485 => x"2d86c72d",
  1486 => x"86c72d86",
  1487 => x"c72d86c7",
  1488 => x"2d86c72d",
  1489 => x"86c72d86",
  1490 => x"c72d86c7",
  1491 => x"2d86c72d",
  1492 => x"86c72d86",
  1493 => x"c72d86c7",
  1494 => x"2d86c72d",
  1495 => x"86c72d86",
  1496 => x"c72d86c7",
  1497 => x"2d86c72d",
  1498 => x"86c72d86",
  1499 => x"c72d86c7",
  1500 => x"2d86c72d",
  1501 => x"86c72d86",
  1502 => x"c72d86c7",
  1503 => x"2d86c72d",
  1504 => x"86c72d86",
  1505 => x"c72d86c7",
  1506 => x"2d86c72d",
  1507 => x"86c72d86",
  1508 => x"c72d86c7",
  1509 => x"2d86c72d",
  1510 => x"86c72d86",
  1511 => x"c72d86c7",
  1512 => x"2d86c72d",
  1513 => x"86c72d86",
  1514 => x"c72d86c7",
  1515 => x"2d86c72d",
  1516 => x"86c72d86",
  1517 => x"c72d86c7",
  1518 => x"2d86c72d",
  1519 => x"86c72d86",
  1520 => x"c72d86c7",
  1521 => x"2d86c72d",
  1522 => x"86c72d86",
  1523 => x"c72d86c7",
  1524 => x"2d86c72d",
  1525 => x"0402dc05",
  1526 => x"0d8059a2",
  1527 => x"902d810b",
  1528 => x"ec0c7a52",
  1529 => x"80e78051",
  1530 => x"80d5e82d",
  1531 => x"80e6e408",
  1532 => x"792e80f7",
  1533 => x"3880e784",
  1534 => x"0870f80c",
  1535 => x"79ff1256",
  1536 => x"59557379",
  1537 => x"2e8b3881",
  1538 => x"1874812a",
  1539 => x"555873f7",
  1540 => x"38f71858",
  1541 => x"81598075",
  1542 => x"2580d038",
  1543 => x"77527351",
  1544 => x"84a82d80",
  1545 => x"e7d85280",
  1546 => x"e7805180",
  1547 => x"d8be2d80",
  1548 => x"e6e40880",
  1549 => x"2e9b3880",
  1550 => x"e7d85783",
  1551 => x"fc567670",
  1552 => x"84055808",
  1553 => x"e80cfc16",
  1554 => x"56758025",
  1555 => x"f138b0d9",
  1556 => x"0480e6e4",
  1557 => x"08598480",
  1558 => x"5580e780",
  1559 => x"5180d88d",
  1560 => x"2dfc8015",
  1561 => x"81155555",
  1562 => x"b0960484",
  1563 => x"0bec0c78",
  1564 => x"802e8e38",
  1565 => x"80e3b451",
  1566 => x"b8e02db6",
  1567 => x"e02db188",
  1568 => x"0480e4b4",
  1569 => x"51b8e02d",
  1570 => x"7880e6e4",
  1571 => x"0c02a405",
  1572 => x"0d0402f0",
  1573 => x"050d840b",
  1574 => x"ec0cb693",
  1575 => x"2db2c12d",
  1576 => x"81f92d83",
  1577 => x"52b5f62d",
  1578 => x"8151858d",
  1579 => x"2dff1252",
  1580 => x"718025f1",
  1581 => x"38840bec",
  1582 => x"0c80e1e4",
  1583 => x"5186a02d",
  1584 => x"80cc882d",
  1585 => x"80e6e408",
  1586 => x"802e80de",
  1587 => x"38afd551",
  1588 => x"80df952d",
  1589 => x"80e3b451",
  1590 => x"b8e02db6",
  1591 => x"cc2db2cd",
  1592 => x"2db8f32d",
  1593 => x"80e3c80b",
  1594 => x"80f52d70",
  1595 => x"842b80e5",
  1596 => x"a0087082",
  1597 => x"2a708106",
  1598 => x"51535654",
  1599 => x"5271802e",
  1600 => x"85387282",
  1601 => x"07537383",
  1602 => x"2a708106",
  1603 => x"51527180",
  1604 => x"2e853872",
  1605 => x"88075372",
  1606 => x"fc0c8652",
  1607 => x"80e6e408",
  1608 => x"83388452",
  1609 => x"71ec0cb1",
  1610 => x"de04800b",
  1611 => x"80e6e40c",
  1612 => x"0290050d",
  1613 => x"0471980c",
  1614 => x"04ffb008",
  1615 => x"80e6e40c",
  1616 => x"04810bff",
  1617 => x"b00c0480",
  1618 => x"0bffb00c",
  1619 => x"0402f405",
  1620 => x"0d80e78c",
  1621 => x"51b4e02d",
  1622 => x"ff0b80e6",
  1623 => x"e4082581",
  1624 => x"883880e6",
  1625 => x"e40881f0",
  1626 => x"2e098106",
  1627 => x"8a38810b",
  1628 => x"80e5980c",
  1629 => x"b3e90480",
  1630 => x"e6e40881",
  1631 => x"e02e0981",
  1632 => x"068a3881",
  1633 => x"0b80e59c",
  1634 => x"0cb3e904",
  1635 => x"80e6e408",
  1636 => x"5280e59c",
  1637 => x"08802e89",
  1638 => x"3880e6e4",
  1639 => x"08818005",
  1640 => x"5271842c",
  1641 => x"728f0653",
  1642 => x"5380e598",
  1643 => x"08802e9a",
  1644 => x"38728429",
  1645 => x"80e4d805",
  1646 => x"72138171",
  1647 => x"2b700973",
  1648 => x"0806730c",
  1649 => x"515353b3",
  1650 => x"dd047284",
  1651 => x"2980e4d8",
  1652 => x"05721383",
  1653 => x"712b7208",
  1654 => x"07720c53",
  1655 => x"53800b80",
  1656 => x"e59c0c80",
  1657 => x"0b80e598",
  1658 => x"0c800b80",
  1659 => x"e6e40c02",
  1660 => x"8c050d04",
  1661 => x"02f8050d",
  1662 => x"80e4d852",
  1663 => x"8f518072",
  1664 => x"70840554",
  1665 => x"0cff1151",
  1666 => x"708025f2",
  1667 => x"38028805",
  1668 => x"0d0402f0",
  1669 => x"050d7551",
  1670 => x"b2c72d70",
  1671 => x"822cfc06",
  1672 => x"80e4d811",
  1673 => x"72109e06",
  1674 => x"71087072",
  1675 => x"2a708306",
  1676 => x"82742b70",
  1677 => x"09740676",
  1678 => x"0c545156",
  1679 => x"57535153",
  1680 => x"b2c12d71",
  1681 => x"80e6e40c",
  1682 => x"0290050d",
  1683 => x"0402fc05",
  1684 => x"0d725180",
  1685 => x"710c800b",
  1686 => x"84120c02",
  1687 => x"84050d04",
  1688 => x"02f0050d",
  1689 => x"75700884",
  1690 => x"12085353",
  1691 => x"53ff5471",
  1692 => x"712ea838",
  1693 => x"b2c72d84",
  1694 => x"13087084",
  1695 => x"29148811",
  1696 => x"70087081",
  1697 => x"ff068418",
  1698 => x"08811187",
  1699 => x"06841a0c",
  1700 => x"53515551",
  1701 => x"5151b2c1",
  1702 => x"2d715473",
  1703 => x"80e6e40c",
  1704 => x"0290050d",
  1705 => x"0402f405",
  1706 => x"0db2c72d",
  1707 => x"e008708b",
  1708 => x"2a708106",
  1709 => x"51525370",
  1710 => x"802ea138",
  1711 => x"80e78c08",
  1712 => x"70842980",
  1713 => x"e7940574",
  1714 => x"81ff0671",
  1715 => x"0c515180",
  1716 => x"e78c0881",
  1717 => x"11870680",
  1718 => x"e78c0c51",
  1719 => x"728c2cbf",
  1720 => x"0680e7b4",
  1721 => x"0c800b80",
  1722 => x"e7b80cb2",
  1723 => x"b92db2c1",
  1724 => x"2d028c05",
  1725 => x"0d0402fc",
  1726 => x"050db2c7",
  1727 => x"2d810b80",
  1728 => x"e7b80cb2",
  1729 => x"c12d80e7",
  1730 => x"b8085170",
  1731 => x"f9380284",
  1732 => x"050d0402",
  1733 => x"fc050d80",
  1734 => x"e78c51b4",
  1735 => x"cd2db3f4",
  1736 => x"2db5a551",
  1737 => x"b2b52d02",
  1738 => x"84050d04",
  1739 => x"02fc050d",
  1740 => x"8fcf5186",
  1741 => x"c72dff11",
  1742 => x"51708025",
  1743 => x"f6380284",
  1744 => x"050d0480",
  1745 => x"e7c40880",
  1746 => x"e6e40c04",
  1747 => x"02fc050d",
  1748 => x"810b80e5",
  1749 => x"a40c8151",
  1750 => x"858d2d02",
  1751 => x"84050d04",
  1752 => x"02fc050d",
  1753 => x"b6ea04b2",
  1754 => x"cd2d8751",
  1755 => x"b4922d80",
  1756 => x"e6e408f3",
  1757 => x"3880e6e4",
  1758 => x"0880e5a4",
  1759 => x"0c80e6e4",
  1760 => x"0851858d",
  1761 => x"2d028405",
  1762 => x"0d0402ec",
  1763 => x"050d7654",
  1764 => x"8052870b",
  1765 => x"881580f5",
  1766 => x"2d565374",
  1767 => x"72248338",
  1768 => x"a0537251",
  1769 => x"83842d81",
  1770 => x"128b1580",
  1771 => x"f52d5452",
  1772 => x"727225de",
  1773 => x"38029405",
  1774 => x"0d0402f0",
  1775 => x"050d80e7",
  1776 => x"c4085481",
  1777 => x"f92d800b",
  1778 => x"80e7c80c",
  1779 => x"7308802e",
  1780 => x"81893882",
  1781 => x"0b80e6f8",
  1782 => x"0c80e7c8",
  1783 => x"088f0680",
  1784 => x"e6f40c73",
  1785 => x"08527183",
  1786 => x"2e963871",
  1787 => x"83268938",
  1788 => x"71812eb0",
  1789 => x"38b8c404",
  1790 => x"71852ea0",
  1791 => x"38b8c404",
  1792 => x"881480f5",
  1793 => x"2d841508",
  1794 => x"80e1fc53",
  1795 => x"545286a0",
  1796 => x"2d718429",
  1797 => x"13700852",
  1798 => x"52b8c804",
  1799 => x"7351b78a",
  1800 => x"2db8c404",
  1801 => x"80e5a008",
  1802 => x"8815082c",
  1803 => x"70810651",
  1804 => x"5271802e",
  1805 => x"883880e2",
  1806 => x"8051b8c1",
  1807 => x"0480e284",
  1808 => x"5186a02d",
  1809 => x"84140851",
  1810 => x"86a02d80",
  1811 => x"e7c80881",
  1812 => x"0580e7c8",
  1813 => x"0c8c1454",
  1814 => x"b7cc0402",
  1815 => x"90050d04",
  1816 => x"7180e7c4",
  1817 => x"0cb7ba2d",
  1818 => x"80e7c808",
  1819 => x"ff0580e7",
  1820 => x"cc0c0402",
  1821 => x"e8050d80",
  1822 => x"e7c40880",
  1823 => x"e7d00857",
  1824 => x"558751b4",
  1825 => x"922d80e6",
  1826 => x"e408812a",
  1827 => x"70810651",
  1828 => x"5271802e",
  1829 => x"a138b99c",
  1830 => x"04b2cd2d",
  1831 => x"8751b492",
  1832 => x"2d80e6e4",
  1833 => x"08f33880",
  1834 => x"e5a40881",
  1835 => x"327080e5",
  1836 => x"a40c5185",
  1837 => x"8d2d80e7",
  1838 => x"b408a006",
  1839 => x"52807225",
  1840 => x"9838b6ac",
  1841 => x"2db2cd2d",
  1842 => x"80e5a408",
  1843 => x"81327080",
  1844 => x"e5a40c70",
  1845 => x"5252858d",
  1846 => x"2d800b80",
  1847 => x"e7bc0c80",
  1848 => x"0b80e7c0",
  1849 => x"0c80e5a4",
  1850 => x"0883ae38",
  1851 => x"80da51b4",
  1852 => x"922d80e6",
  1853 => x"e408802e",
  1854 => x"8c3880e7",
  1855 => x"bc088180",
  1856 => x"0780e7bc",
  1857 => x"0c80d951",
  1858 => x"b4922d80",
  1859 => x"e6e40880",
  1860 => x"2e8c3880",
  1861 => x"e7bc0880",
  1862 => x"c00780e7",
  1863 => x"bc0c8194",
  1864 => x"51b4922d",
  1865 => x"80e6e408",
  1866 => x"802e8b38",
  1867 => x"80e7bc08",
  1868 => x"900780e7",
  1869 => x"bc0c8191",
  1870 => x"51b4922d",
  1871 => x"80e6e408",
  1872 => x"802e8b38",
  1873 => x"80e7bc08",
  1874 => x"a00780e7",
  1875 => x"bc0c81f5",
  1876 => x"51b4922d",
  1877 => x"80e6e408",
  1878 => x"802e8b38",
  1879 => x"80e7bc08",
  1880 => x"810780e7",
  1881 => x"bc0c81f2",
  1882 => x"51b4922d",
  1883 => x"80e6e408",
  1884 => x"802e8b38",
  1885 => x"80e7bc08",
  1886 => x"820780e7",
  1887 => x"bc0c81eb",
  1888 => x"51b4922d",
  1889 => x"80e6e408",
  1890 => x"802e8b38",
  1891 => x"80e7bc08",
  1892 => x"840780e7",
  1893 => x"bc0c81f4",
  1894 => x"51b4922d",
  1895 => x"80e6e408",
  1896 => x"802e8b38",
  1897 => x"80e7bc08",
  1898 => x"880780e7",
  1899 => x"bc0c80d8",
  1900 => x"51b4922d",
  1901 => x"80e6e408",
  1902 => x"802e8c38",
  1903 => x"80e7c008",
  1904 => x"81800780",
  1905 => x"e7c00c92",
  1906 => x"51b4922d",
  1907 => x"80e6e408",
  1908 => x"802e8c38",
  1909 => x"80e7c008",
  1910 => x"80c00780",
  1911 => x"e7c00c94",
  1912 => x"51b4922d",
  1913 => x"80e6e408",
  1914 => x"802e8b38",
  1915 => x"80e7c008",
  1916 => x"900780e7",
  1917 => x"c00c9151",
  1918 => x"b4922d80",
  1919 => x"e6e40880",
  1920 => x"2e8b3880",
  1921 => x"e7c008a0",
  1922 => x"0780e7c0",
  1923 => x"0c9d51b4",
  1924 => x"922d80e6",
  1925 => x"e408802e",
  1926 => x"8b3880e7",
  1927 => x"c0088107",
  1928 => x"80e7c00c",
  1929 => x"9b51b492",
  1930 => x"2d80e6e4",
  1931 => x"08802e8b",
  1932 => x"3880e7c0",
  1933 => x"08820780",
  1934 => x"e7c00c9c",
  1935 => x"51b4922d",
  1936 => x"80e6e408",
  1937 => x"802e8b38",
  1938 => x"80e7c008",
  1939 => x"840780e7",
  1940 => x"c00ca351",
  1941 => x"b4922d80",
  1942 => x"e6e40880",
  1943 => x"2e8b3880",
  1944 => x"e7c00888",
  1945 => x"0780e7c0",
  1946 => x"0c9651b4",
  1947 => x"922d80e6",
  1948 => x"e408802e",
  1949 => x"843894bf",
  1950 => x"2d9e51b4",
  1951 => x"922d80e6",
  1952 => x"e408802e",
  1953 => x"843886ee",
  1954 => x"2d81fd51",
  1955 => x"b4922d81",
  1956 => x"fa51b492",
  1957 => x"2d80c3c1",
  1958 => x"0481f551",
  1959 => x"b4922d80",
  1960 => x"e6e40881",
  1961 => x"2a708106",
  1962 => x"5152718e",
  1963 => x"3880e7b4",
  1964 => x"08900652",
  1965 => x"80722580",
  1966 => x"c23880e7",
  1967 => x"b4089006",
  1968 => x"52807225",
  1969 => x"8438b6ac",
  1970 => x"2d80e7cc",
  1971 => x"08527180",
  1972 => x"2e8a38ff",
  1973 => x"1280e7cc",
  1974 => x"0cbdfb04",
  1975 => x"80e7c808",
  1976 => x"1080e7c8",
  1977 => x"08057084",
  1978 => x"29165152",
  1979 => x"88120880",
  1980 => x"2e8938ff",
  1981 => x"51881208",
  1982 => x"52712d81",
  1983 => x"f251b492",
  1984 => x"2d80e6e4",
  1985 => x"08812a70",
  1986 => x"81065152",
  1987 => x"718e3880",
  1988 => x"e7b40888",
  1989 => x"06528072",
  1990 => x"2580c338",
  1991 => x"80e7b408",
  1992 => x"88065280",
  1993 => x"72258438",
  1994 => x"b6ac2d80",
  1995 => x"e7c808ff",
  1996 => x"1180e7cc",
  1997 => x"08565353",
  1998 => x"7372258a",
  1999 => x"38811480",
  2000 => x"e7cc0cbe",
  2001 => x"de047210",
  2002 => x"13708429",
  2003 => x"16515288",
  2004 => x"1208802e",
  2005 => x"8938fe51",
  2006 => x"88120852",
  2007 => x"712d81fd",
  2008 => x"51b4922d",
  2009 => x"80e6e408",
  2010 => x"812a7081",
  2011 => x"06515271",
  2012 => x"802eb138",
  2013 => x"80e7cc08",
  2014 => x"802e8a38",
  2015 => x"800b80e7",
  2016 => x"cc0cbfa4",
  2017 => x"0480e7c8",
  2018 => x"081080e7",
  2019 => x"c8080570",
  2020 => x"84291651",
  2021 => x"52881208",
  2022 => x"802e8938",
  2023 => x"fd518812",
  2024 => x"0852712d",
  2025 => x"81fa51b4",
  2026 => x"922d80e6",
  2027 => x"e408812a",
  2028 => x"70810651",
  2029 => x"5271802e",
  2030 => x"b13880e7",
  2031 => x"c808ff11",
  2032 => x"545280e7",
  2033 => x"cc087325",
  2034 => x"89387280",
  2035 => x"e7cc0cbf",
  2036 => x"ea047110",
  2037 => x"12708429",
  2038 => x"16515288",
  2039 => x"1208802e",
  2040 => x"8938fc51",
  2041 => x"88120852",
  2042 => x"712d80e7",
  2043 => x"cc087053",
  2044 => x"5473802e",
  2045 => x"8a388c15",
  2046 => x"ff155555",
  2047 => x"bff10482",
  2048 => x"0b80e6f8",
  2049 => x"0c718f06",
  2050 => x"80e6f40c",
  2051 => x"81eb51b4",
  2052 => x"922d80e6",
  2053 => x"e408812a",
  2054 => x"70810651",
  2055 => x"5271802e",
  2056 => x"ad387408",
  2057 => x"852e0981",
  2058 => x"06a43888",
  2059 => x"1580f52d",
  2060 => x"ff055271",
  2061 => x"881681b7",
  2062 => x"2d71982b",
  2063 => x"52718025",
  2064 => x"8838800b",
  2065 => x"881681b7",
  2066 => x"2d7451b7",
  2067 => x"8a2d81f4",
  2068 => x"51b4922d",
  2069 => x"80e6e408",
  2070 => x"812a7081",
  2071 => x"06515271",
  2072 => x"802eb338",
  2073 => x"7408852e",
  2074 => x"098106aa",
  2075 => x"38881580",
  2076 => x"f52d8105",
  2077 => x"52718816",
  2078 => x"81b72d71",
  2079 => x"81ff068b",
  2080 => x"1680f52d",
  2081 => x"54527272",
  2082 => x"27873872",
  2083 => x"881681b7",
  2084 => x"2d7451b7",
  2085 => x"8a2d80da",
  2086 => x"51b4922d",
  2087 => x"80e6e408",
  2088 => x"812a7081",
  2089 => x"06515271",
  2090 => x"8e3880e7",
  2091 => x"b4088106",
  2092 => x"52807225",
  2093 => x"81c23880",
  2094 => x"e7c40880",
  2095 => x"e7b40881",
  2096 => x"06535380",
  2097 => x"72258438",
  2098 => x"b6ac2d80",
  2099 => x"e7cc0854",
  2100 => x"73802e8b",
  2101 => x"388c13ff",
  2102 => x"15555380",
  2103 => x"c1d00472",
  2104 => x"08527182",
  2105 => x"2ea83871",
  2106 => x"82268a38",
  2107 => x"71812ead",
  2108 => x"3880c2f8",
  2109 => x"0471832e",
  2110 => x"b7387184",
  2111 => x"2e098106",
  2112 => x"80f63888",
  2113 => x"130851b8",
  2114 => x"e02d80c2",
  2115 => x"f80480e7",
  2116 => x"cc085188",
  2117 => x"13085271",
  2118 => x"2d80c2f8",
  2119 => x"04810b88",
  2120 => x"14082b80",
  2121 => x"e5a00832",
  2122 => x"80e5a00c",
  2123 => x"80c2cb04",
  2124 => x"881380f5",
  2125 => x"2d81058b",
  2126 => x"1480f52d",
  2127 => x"53547174",
  2128 => x"24833880",
  2129 => x"54738814",
  2130 => x"81b72db7",
  2131 => x"ba2d80c2",
  2132 => x"f8047508",
  2133 => x"802ea438",
  2134 => x"750851b4",
  2135 => x"922d80e6",
  2136 => x"e4088106",
  2137 => x"5271802e",
  2138 => x"8c3880e7",
  2139 => x"cc085184",
  2140 => x"16085271",
  2141 => x"2d881656",
  2142 => x"75d83880",
  2143 => x"54800b80",
  2144 => x"e6f80c73",
  2145 => x"8f0680e6",
  2146 => x"f40ca052",
  2147 => x"7380e7cc",
  2148 => x"082e0981",
  2149 => x"06993880",
  2150 => x"e7c808ff",
  2151 => x"05743270",
  2152 => x"09810570",
  2153 => x"72079f2a",
  2154 => x"91713151",
  2155 => x"51535371",
  2156 => x"5183842d",
  2157 => x"8114548e",
  2158 => x"7425c238",
  2159 => x"80e5a408",
  2160 => x"527180e6",
  2161 => x"e40c0298",
  2162 => x"050d0402",
  2163 => x"f4050dd4",
  2164 => x"5281ff72",
  2165 => x"0c710853",
  2166 => x"81ff720c",
  2167 => x"72882b83",
  2168 => x"fe800672",
  2169 => x"087081ff",
  2170 => x"06515253",
  2171 => x"81ff720c",
  2172 => x"72710788",
  2173 => x"2b720870",
  2174 => x"81ff0651",
  2175 => x"525381ff",
  2176 => x"720c7271",
  2177 => x"07882b72",
  2178 => x"087081ff",
  2179 => x"06720780",
  2180 => x"e6e40c52",
  2181 => x"53028c05",
  2182 => x"0d0402f4",
  2183 => x"050d7476",
  2184 => x"7181ff06",
  2185 => x"d40c5353",
  2186 => x"80e7d408",
  2187 => x"85387189",
  2188 => x"2b527198",
  2189 => x"2ad40c71",
  2190 => x"902a7081",
  2191 => x"ff06d40c",
  2192 => x"5171882a",
  2193 => x"7081ff06",
  2194 => x"d40c5171",
  2195 => x"81ff06d4",
  2196 => x"0c72902a",
  2197 => x"7081ff06",
  2198 => x"d40c51d4",
  2199 => x"087081ff",
  2200 => x"06515182",
  2201 => x"b8bf5270",
  2202 => x"81ff2e09",
  2203 => x"81069438",
  2204 => x"81ff0bd4",
  2205 => x"0cd40870",
  2206 => x"81ff06ff",
  2207 => x"14545151",
  2208 => x"71e53870",
  2209 => x"80e6e40c",
  2210 => x"028c050d",
  2211 => x"0402fc05",
  2212 => x"0d81c751",
  2213 => x"81ff0bd4",
  2214 => x"0cff1151",
  2215 => x"708025f4",
  2216 => x"38028405",
  2217 => x"0d0402f4",
  2218 => x"050d81ff",
  2219 => x"0bd40c93",
  2220 => x"53805287",
  2221 => x"fc80c151",
  2222 => x"80c49a2d",
  2223 => x"80e6e408",
  2224 => x"8c3881ff",
  2225 => x"0bd40c81",
  2226 => x"5380c5d7",
  2227 => x"0480c58d",
  2228 => x"2dff1353",
  2229 => x"72db3872",
  2230 => x"80e6e40c",
  2231 => x"028c050d",
  2232 => x"0402ec05",
  2233 => x"0d810b80",
  2234 => x"e7d40c84",
  2235 => x"54d00870",
  2236 => x"8f2a7081",
  2237 => x"06515153",
  2238 => x"72f33872",
  2239 => x"d00c80c5",
  2240 => x"8d2d80e2",
  2241 => x"885186a0",
  2242 => x"2dd00870",
  2243 => x"8f2a7081",
  2244 => x"06515153",
  2245 => x"72f33881",
  2246 => x"0bd00cb1",
  2247 => x"53805284",
  2248 => x"d480c051",
  2249 => x"80c49a2d",
  2250 => x"80e6e408",
  2251 => x"812e9438",
  2252 => x"72822e80",
  2253 => x"c438ff13",
  2254 => x"5372e238",
  2255 => x"ff145473",
  2256 => x"ffab3880",
  2257 => x"c58d2d83",
  2258 => x"aa52849c",
  2259 => x"80c85180",
  2260 => x"c49a2d80",
  2261 => x"e6e40881",
  2262 => x"2e098106",
  2263 => x"943880c3",
  2264 => x"cb2d80e6",
  2265 => x"e40883ff",
  2266 => x"ff065372",
  2267 => x"83aa2ea3",
  2268 => x"3880c5a6",
  2269 => x"2d80c78d",
  2270 => x"0480e294",
  2271 => x"5186a02d",
  2272 => x"805380c8",
  2273 => x"eb0480e2",
  2274 => x"ac5186a0",
  2275 => x"2d805480",
  2276 => x"c8bb0481",
  2277 => x"ff0bd40c",
  2278 => x"b15480c5",
  2279 => x"8d2d8fcf",
  2280 => x"53805287",
  2281 => x"fc80f751",
  2282 => x"80c49a2d",
  2283 => x"80e6e408",
  2284 => x"5580e6e4",
  2285 => x"08812e09",
  2286 => x"81069e38",
  2287 => x"81ff0bd4",
  2288 => x"0c820a52",
  2289 => x"849c80e9",
  2290 => x"5180c49a",
  2291 => x"2d80e6e4",
  2292 => x"08802e8f",
  2293 => x"3880c58d",
  2294 => x"2dff1353",
  2295 => x"72c33880",
  2296 => x"c8ae0481",
  2297 => x"ff0bd40c",
  2298 => x"80e6e408",
  2299 => x"5287fc80",
  2300 => x"fa5180c4",
  2301 => x"9a2d80e6",
  2302 => x"e408b338",
  2303 => x"81ff0bd4",
  2304 => x"0cd40853",
  2305 => x"81ff0bd4",
  2306 => x"0c81ff0b",
  2307 => x"d40c81ff",
  2308 => x"0bd40c81",
  2309 => x"ff0bd40c",
  2310 => x"72862a70",
  2311 => x"81067656",
  2312 => x"51537297",
  2313 => x"3880e6e4",
  2314 => x"085480c8",
  2315 => x"bb047382",
  2316 => x"2efed338",
  2317 => x"ff145473",
  2318 => x"fee03873",
  2319 => x"80e7d40c",
  2320 => x"738c3881",
  2321 => x"5287fc80",
  2322 => x"d05180c4",
  2323 => x"9a2d81ff",
  2324 => x"0bd40cd0",
  2325 => x"08708f2a",
  2326 => x"70810651",
  2327 => x"515372f3",
  2328 => x"3872d00c",
  2329 => x"81ff0bd4",
  2330 => x"0c815372",
  2331 => x"80e6e40c",
  2332 => x"0294050d",
  2333 => x"0402e805",
  2334 => x"0d785580",
  2335 => x"5681ff0b",
  2336 => x"d40cd008",
  2337 => x"708f2a70",
  2338 => x"81065151",
  2339 => x"5372f338",
  2340 => x"82810bd0",
  2341 => x"0c81ff0b",
  2342 => x"d40c7752",
  2343 => x"87fc80d1",
  2344 => x"5180c49a",
  2345 => x"2d80dbc6",
  2346 => x"df5480e6",
  2347 => x"e408802e",
  2348 => x"8c3880e2",
  2349 => x"cc5186a0",
  2350 => x"2d80ca93",
  2351 => x"0481ff0b",
  2352 => x"d40cd408",
  2353 => x"7081ff06",
  2354 => x"51537281",
  2355 => x"fe2e0981",
  2356 => x"06a03880",
  2357 => x"ff5380c3",
  2358 => x"cb2d80e6",
  2359 => x"e4087570",
  2360 => x"8405570c",
  2361 => x"ff135372",
  2362 => x"8025eb38",
  2363 => x"815680c9",
  2364 => x"f804ff14",
  2365 => x"5473c638",
  2366 => x"81ff0bd4",
  2367 => x"0c81ff0b",
  2368 => x"d40cd008",
  2369 => x"708f2a70",
  2370 => x"81065151",
  2371 => x"5372f338",
  2372 => x"72d00c75",
  2373 => x"80e6e40c",
  2374 => x"0298050d",
  2375 => x"0402e805",
  2376 => x"0d77797b",
  2377 => x"58555580",
  2378 => x"53727625",
  2379 => x"a5387470",
  2380 => x"81055680",
  2381 => x"f52d7470",
  2382 => x"81055680",
  2383 => x"f52d5252",
  2384 => x"71712e87",
  2385 => x"38815180",
  2386 => x"cad40481",
  2387 => x"135380ca",
  2388 => x"a9048051",
  2389 => x"7080e6e4",
  2390 => x"0c029805",
  2391 => x"0d0402ec",
  2392 => x"050d7655",
  2393 => x"74802e80",
  2394 => x"c4389a15",
  2395 => x"80e02d51",
  2396 => x"80d9992d",
  2397 => x"80e6e408",
  2398 => x"80e6e408",
  2399 => x"80ee880c",
  2400 => x"80e6e408",
  2401 => x"545480ed",
  2402 => x"e408802e",
  2403 => x"9b389415",
  2404 => x"80e02d51",
  2405 => x"80d9992d",
  2406 => x"80e6e408",
  2407 => x"902b83ff",
  2408 => x"f00a0670",
  2409 => x"75075153",
  2410 => x"7280ee88",
  2411 => x"0c80ee88",
  2412 => x"08537280",
  2413 => x"2e9e3880",
  2414 => x"eddc08fe",
  2415 => x"14712980",
  2416 => x"edf00805",
  2417 => x"80ee8c0c",
  2418 => x"70842b80",
  2419 => x"ede80c54",
  2420 => x"80cc8304",
  2421 => x"80edf408",
  2422 => x"80ee880c",
  2423 => x"80edf808",
  2424 => x"80ee8c0c",
  2425 => x"80ede408",
  2426 => x"802e8c38",
  2427 => x"80eddc08",
  2428 => x"842b5380",
  2429 => x"cbfe0480",
  2430 => x"edfc0884",
  2431 => x"2b537280",
  2432 => x"ede80c02",
  2433 => x"94050d04",
  2434 => x"02d8050d",
  2435 => x"800b80ed",
  2436 => x"e40c8454",
  2437 => x"80c5e12d",
  2438 => x"80e6e408",
  2439 => x"802e9938",
  2440 => x"80e7d852",
  2441 => x"805180c8",
  2442 => x"f52d80e6",
  2443 => x"e408802e",
  2444 => x"8738fe54",
  2445 => x"80ccc004",
  2446 => x"ff145473",
  2447 => x"8024d538",
  2448 => x"738e3880",
  2449 => x"e2dc5186",
  2450 => x"a02d7355",
  2451 => x"80d2a404",
  2452 => x"8056810b",
  2453 => x"80ee900c",
  2454 => x"885380e2",
  2455 => x"f05280e8",
  2456 => x"8e5180ca",
  2457 => x"9d2d80e6",
  2458 => x"e408762e",
  2459 => x"09810689",
  2460 => x"3880e6e4",
  2461 => x"0880ee90",
  2462 => x"0c885380",
  2463 => x"e2fc5280",
  2464 => x"e8aa5180",
  2465 => x"ca9d2d80",
  2466 => x"e6e40889",
  2467 => x"3880e6e4",
  2468 => x"0880ee90",
  2469 => x"0c80ee90",
  2470 => x"08802e81",
  2471 => x"853880eb",
  2472 => x"9e0b80f5",
  2473 => x"2d80eb9f",
  2474 => x"0b80f52d",
  2475 => x"71982b71",
  2476 => x"902b0780",
  2477 => x"eba00b80",
  2478 => x"f52d7088",
  2479 => x"2b720780",
  2480 => x"eba10b80",
  2481 => x"f52d7107",
  2482 => x"80ebd60b",
  2483 => x"80f52d80",
  2484 => x"ebd70b80",
  2485 => x"f52d7188",
  2486 => x"2b07535f",
  2487 => x"54525a56",
  2488 => x"57557381",
  2489 => x"abaa2e09",
  2490 => x"81069038",
  2491 => x"755180d8",
  2492 => x"e82d80e6",
  2493 => x"e4085680",
  2494 => x"ce8a0473",
  2495 => x"82d4d52e",
  2496 => x"893880e3",
  2497 => x"885180ce",
  2498 => x"da0480e7",
  2499 => x"d8527551",
  2500 => x"80c8f52d",
  2501 => x"80e6e408",
  2502 => x"5580e6e4",
  2503 => x"08802e84",
  2504 => x"83388853",
  2505 => x"80e2fc52",
  2506 => x"80e8aa51",
  2507 => x"80ca9d2d",
  2508 => x"80e6e408",
  2509 => x"8b38810b",
  2510 => x"80ede40c",
  2511 => x"80cee104",
  2512 => x"885380e2",
  2513 => x"f05280e8",
  2514 => x"8e5180ca",
  2515 => x"9d2d80e6",
  2516 => x"e408802e",
  2517 => x"8c3880e3",
  2518 => x"9c5186a0",
  2519 => x"2d80cfc0",
  2520 => x"0480ebd6",
  2521 => x"0b80f52d",
  2522 => x"547380d5",
  2523 => x"2e098106",
  2524 => x"80ce3880",
  2525 => x"ebd70b80",
  2526 => x"f52d5473",
  2527 => x"81aa2e09",
  2528 => x"8106bd38",
  2529 => x"800b80e7",
  2530 => x"d80b80f5",
  2531 => x"2d565474",
  2532 => x"81e92e83",
  2533 => x"38815474",
  2534 => x"81eb2e8c",
  2535 => x"38805573",
  2536 => x"752e0981",
  2537 => x"0682fd38",
  2538 => x"80e7e30b",
  2539 => x"80f52d55",
  2540 => x"748e3880",
  2541 => x"e7e40b80",
  2542 => x"f52d5473",
  2543 => x"822e8738",
  2544 => x"805580d2",
  2545 => x"a40480e7",
  2546 => x"e50b80f5",
  2547 => x"2d7080ed",
  2548 => x"dc0cff05",
  2549 => x"80ede00c",
  2550 => x"80e7e60b",
  2551 => x"80f52d80",
  2552 => x"e7e70b80",
  2553 => x"f52d5876",
  2554 => x"05778280",
  2555 => x"29057080",
  2556 => x"edec0c80",
  2557 => x"e7e80b80",
  2558 => x"f52d7080",
  2559 => x"ee800c80",
  2560 => x"ede40859",
  2561 => x"57587680",
  2562 => x"2e81b938",
  2563 => x"885380e2",
  2564 => x"fc5280e8",
  2565 => x"aa5180ca",
  2566 => x"9d2d80e6",
  2567 => x"e4088284",
  2568 => x"3880eddc",
  2569 => x"0870842b",
  2570 => x"80ede80c",
  2571 => x"7080edfc",
  2572 => x"0c80e7fd",
  2573 => x"0b80f52d",
  2574 => x"80e7fc0b",
  2575 => x"80f52d71",
  2576 => x"82802905",
  2577 => x"80e7fe0b",
  2578 => x"80f52d70",
  2579 => x"84808029",
  2580 => x"1280e7ff",
  2581 => x"0b80f52d",
  2582 => x"7081800a",
  2583 => x"29127080",
  2584 => x"ee840c80",
  2585 => x"ee800871",
  2586 => x"2980edec",
  2587 => x"08057080",
  2588 => x"edf00c80",
  2589 => x"e8850b80",
  2590 => x"f52d80e8",
  2591 => x"840b80f5",
  2592 => x"2d718280",
  2593 => x"290580e8",
  2594 => x"860b80f5",
  2595 => x"2d708480",
  2596 => x"80291280",
  2597 => x"e8870b80",
  2598 => x"f52d7098",
  2599 => x"2b81f00a",
  2600 => x"06720570",
  2601 => x"80edf40c",
  2602 => x"fe117e29",
  2603 => x"770580ed",
  2604 => x"f80c5259",
  2605 => x"5243545e",
  2606 => x"51525952",
  2607 => x"5d575957",
  2608 => x"80d29c04",
  2609 => x"80e7ea0b",
  2610 => x"80f52d80",
  2611 => x"e7e90b80",
  2612 => x"f52d7182",
  2613 => x"80290570",
  2614 => x"80ede80c",
  2615 => x"70a02983",
  2616 => x"ff057089",
  2617 => x"2a7080ed",
  2618 => x"fc0c80e7",
  2619 => x"ef0b80f5",
  2620 => x"2d80e7ee",
  2621 => x"0b80f52d",
  2622 => x"71828029",
  2623 => x"057080ee",
  2624 => x"840c7b71",
  2625 => x"291e7080",
  2626 => x"edf80c7d",
  2627 => x"80edf40c",
  2628 => x"730580ed",
  2629 => x"f00c555e",
  2630 => x"51515555",
  2631 => x"805180ca",
  2632 => x"de2d8155",
  2633 => x"7480e6e4",
  2634 => x"0c02a805",
  2635 => x"0d0402ec",
  2636 => x"050d7670",
  2637 => x"872c7180",
  2638 => x"ff065556",
  2639 => x"5480ede4",
  2640 => x"088a3873",
  2641 => x"882c7481",
  2642 => x"ff065455",
  2643 => x"80e7d852",
  2644 => x"80edec08",
  2645 => x"155180c8",
  2646 => x"f52d80e6",
  2647 => x"e4085480",
  2648 => x"e6e40880",
  2649 => x"2ebb3880",
  2650 => x"ede40880",
  2651 => x"2e9c3872",
  2652 => x"842980e7",
  2653 => x"d8057008",
  2654 => x"525380d8",
  2655 => x"e82d80e6",
  2656 => x"e408f00a",
  2657 => x"065380d3",
  2658 => x"9f047210",
  2659 => x"80e7d805",
  2660 => x"7080e02d",
  2661 => x"525380d9",
  2662 => x"992d80e6",
  2663 => x"e4085372",
  2664 => x"547380e6",
  2665 => x"e40c0294",
  2666 => x"050d0402",
  2667 => x"e0050d79",
  2668 => x"70842c80",
  2669 => x"ee8c0805",
  2670 => x"718f0652",
  2671 => x"5553728b",
  2672 => x"3880e7d8",
  2673 => x"52735180",
  2674 => x"c8f52d72",
  2675 => x"a02980e7",
  2676 => x"d8055480",
  2677 => x"7480f52d",
  2678 => x"56537473",
  2679 => x"2e833881",
  2680 => x"537481e5",
  2681 => x"2e81f538",
  2682 => x"81707406",
  2683 => x"54587280",
  2684 => x"2e81e938",
  2685 => x"8b1480f5",
  2686 => x"2d70832a",
  2687 => x"79065856",
  2688 => x"769c3880",
  2689 => x"e5a80853",
  2690 => x"72893872",
  2691 => x"80ebd80b",
  2692 => x"81b72d76",
  2693 => x"80e5a80c",
  2694 => x"735380d5",
  2695 => x"de04758f",
  2696 => x"2e098106",
  2697 => x"81b63874",
  2698 => x"9f068d29",
  2699 => x"80ebcb11",
  2700 => x"51538114",
  2701 => x"80f52d73",
  2702 => x"70810555",
  2703 => x"81b72d83",
  2704 => x"1480f52d",
  2705 => x"73708105",
  2706 => x"5581b72d",
  2707 => x"851480f5",
  2708 => x"2d737081",
  2709 => x"055581b7",
  2710 => x"2d871480",
  2711 => x"f52d7370",
  2712 => x"81055581",
  2713 => x"b72d8914",
  2714 => x"80f52d73",
  2715 => x"70810555",
  2716 => x"81b72d8e",
  2717 => x"1480f52d",
  2718 => x"73708105",
  2719 => x"5581b72d",
  2720 => x"901480f5",
  2721 => x"2d737081",
  2722 => x"055581b7",
  2723 => x"2d921480",
  2724 => x"f52d7370",
  2725 => x"81055581",
  2726 => x"b72d9414",
  2727 => x"80f52d73",
  2728 => x"70810555",
  2729 => x"81b72d96",
  2730 => x"1480f52d",
  2731 => x"73708105",
  2732 => x"5581b72d",
  2733 => x"981480f5",
  2734 => x"2d737081",
  2735 => x"055581b7",
  2736 => x"2d9c1480",
  2737 => x"f52d7370",
  2738 => x"81055581",
  2739 => x"b72d9e14",
  2740 => x"80f52d73",
  2741 => x"81b72d77",
  2742 => x"80e5a80c",
  2743 => x"80537280",
  2744 => x"e6e40c02",
  2745 => x"a0050d04",
  2746 => x"02cc050d",
  2747 => x"7e605e5a",
  2748 => x"800b80ee",
  2749 => x"880880ee",
  2750 => x"8c08595c",
  2751 => x"56805880",
  2752 => x"ede80878",
  2753 => x"2e81be38",
  2754 => x"778f06a0",
  2755 => x"17575473",
  2756 => x"923880e7",
  2757 => x"d8527651",
  2758 => x"81175780",
  2759 => x"c8f52d80",
  2760 => x"e7d85680",
  2761 => x"7680f52d",
  2762 => x"56547474",
  2763 => x"2e833881",
  2764 => x"547481e5",
  2765 => x"2e818238",
  2766 => x"81707506",
  2767 => x"555c7380",
  2768 => x"2e80f638",
  2769 => x"8b1680f5",
  2770 => x"2d980659",
  2771 => x"7880ea38",
  2772 => x"8b537c52",
  2773 => x"755180ca",
  2774 => x"9d2d80e6",
  2775 => x"e40880d9",
  2776 => x"389c1608",
  2777 => x"5180d8e8",
  2778 => x"2d80e6e4",
  2779 => x"08841b0c",
  2780 => x"9a1680e0",
  2781 => x"2d5180d9",
  2782 => x"992d80e6",
  2783 => x"e40880e6",
  2784 => x"e408881c",
  2785 => x"0c80e6e4",
  2786 => x"08555580",
  2787 => x"ede40880",
  2788 => x"2e9a3894",
  2789 => x"1680e02d",
  2790 => x"5180d999",
  2791 => x"2d80e6e4",
  2792 => x"08902b83",
  2793 => x"fff00a06",
  2794 => x"70165154",
  2795 => x"73881b0c",
  2796 => x"787a0c7b",
  2797 => x"5480d883",
  2798 => x"04811858",
  2799 => x"80ede808",
  2800 => x"7826fec4",
  2801 => x"3880ede4",
  2802 => x"08802eb5",
  2803 => x"387a5180",
  2804 => x"d2ae2d80",
  2805 => x"e6e40880",
  2806 => x"e6e40880",
  2807 => x"fffffff8",
  2808 => x"06555b73",
  2809 => x"80ffffff",
  2810 => x"f82e9638",
  2811 => x"80e6e408",
  2812 => x"fe0580ed",
  2813 => x"dc082980",
  2814 => x"edf00805",
  2815 => x"5780d5fd",
  2816 => x"04805473",
  2817 => x"80e6e40c",
  2818 => x"02b4050d",
  2819 => x"0402f405",
  2820 => x"0d747008",
  2821 => x"8105710c",
  2822 => x"700880ed",
  2823 => x"e0080653",
  2824 => x"53719038",
  2825 => x"88130851",
  2826 => x"80d2ae2d",
  2827 => x"80e6e408",
  2828 => x"88140c81",
  2829 => x"0b80e6e4",
  2830 => x"0c028c05",
  2831 => x"0d0402f0",
  2832 => x"050d7588",
  2833 => x"1108fe05",
  2834 => x"80eddc08",
  2835 => x"2980edf0",
  2836 => x"08117208",
  2837 => x"80ede008",
  2838 => x"06057955",
  2839 => x"53545480",
  2840 => x"c8f52d02",
  2841 => x"90050d04",
  2842 => x"02f4050d",
  2843 => x"7470882a",
  2844 => x"83fe8006",
  2845 => x"7072982a",
  2846 => x"0772882b",
  2847 => x"87fc8080",
  2848 => x"0673982b",
  2849 => x"81f00a06",
  2850 => x"71730707",
  2851 => x"80e6e40c",
  2852 => x"56515351",
  2853 => x"028c050d",
  2854 => x"0402f805",
  2855 => x"0d028e05",
  2856 => x"80f52d74",
  2857 => x"882b0770",
  2858 => x"83ffff06",
  2859 => x"80e6e40c",
  2860 => x"51028805",
  2861 => x"0d0402f4",
  2862 => x"050d7476",
  2863 => x"78535452",
  2864 => x"80712597",
  2865 => x"38727081",
  2866 => x"055480f5",
  2867 => x"2d727081",
  2868 => x"055481b7",
  2869 => x"2dff1151",
  2870 => x"70eb3880",
  2871 => x"7281b72d",
  2872 => x"028c050d",
  2873 => x"0402e805",
  2874 => x"0d775680",
  2875 => x"70565473",
  2876 => x"7624b738",
  2877 => x"80ede808",
  2878 => x"742eaf38",
  2879 => x"735180d3",
  2880 => x"ab2d80e6",
  2881 => x"e40880e6",
  2882 => x"e4080981",
  2883 => x"057080e6",
  2884 => x"e408079f",
  2885 => x"2a770581",
  2886 => x"17575753",
  2887 => x"53747624",
  2888 => x"893880ed",
  2889 => x"e8087426",
  2890 => x"d3387280",
  2891 => x"e6e40c02",
  2892 => x"98050d04",
  2893 => x"02f0050d",
  2894 => x"80e6e008",
  2895 => x"165180d9",
  2896 => x"e52d80e6",
  2897 => x"e408802e",
  2898 => x"a0388b53",
  2899 => x"80e6e408",
  2900 => x"5280ebd8",
  2901 => x"5180d9b6",
  2902 => x"2d80ee94",
  2903 => x"08547380",
  2904 => x"2e873880",
  2905 => x"ebd85173",
  2906 => x"2d029005",
  2907 => x"0d0402dc",
  2908 => x"050d8070",
  2909 => x"5a557480",
  2910 => x"e6e00825",
  2911 => x"b53880ed",
  2912 => x"e808752e",
  2913 => x"ad387851",
  2914 => x"80d3ab2d",
  2915 => x"80e6e408",
  2916 => x"09810570",
  2917 => x"80e6e408",
  2918 => x"079f2a76",
  2919 => x"05811b5b",
  2920 => x"56547480",
  2921 => x"e6e00825",
  2922 => x"893880ed",
  2923 => x"e8087926",
  2924 => x"d5388055",
  2925 => x"7880ede8",
  2926 => x"082781e4",
  2927 => x"38785180",
  2928 => x"d3ab2d80",
  2929 => x"e6e40880",
  2930 => x"2e81b438",
  2931 => x"80e6e408",
  2932 => x"8b0580f5",
  2933 => x"2d70842a",
  2934 => x"70810677",
  2935 => x"1078842b",
  2936 => x"80ebd80b",
  2937 => x"80f52d5c",
  2938 => x"5c535155",
  2939 => x"5673802e",
  2940 => x"80ce3874",
  2941 => x"16822b80",
  2942 => x"ddc40b80",
  2943 => x"e5b4120c",
  2944 => x"54777531",
  2945 => x"1080ee98",
  2946 => x"11555690",
  2947 => x"74708105",
  2948 => x"5681b72d",
  2949 => x"a07481b7",
  2950 => x"2d7681ff",
  2951 => x"06811658",
  2952 => x"5473802e",
  2953 => x"8b389c53",
  2954 => x"80ebd852",
  2955 => x"80dcb704",
  2956 => x"8b5380e6",
  2957 => x"e4085280",
  2958 => x"ee9a1651",
  2959 => x"80dcf504",
  2960 => x"7416822b",
  2961 => x"80dab40b",
  2962 => x"80e5b412",
  2963 => x"0c547681",
  2964 => x"ff068116",
  2965 => x"58547380",
  2966 => x"2e8b389c",
  2967 => x"5380ebd8",
  2968 => x"5280dcec",
  2969 => x"048b5380",
  2970 => x"e6e40852",
  2971 => x"77753110",
  2972 => x"80ee9805",
  2973 => x"51765580",
  2974 => x"d9b62d80",
  2975 => x"dd940474",
  2976 => x"90297531",
  2977 => x"701080ee",
  2978 => x"98055154",
  2979 => x"80e6e408",
  2980 => x"7481b72d",
  2981 => x"81195974",
  2982 => x"8b24a438",
  2983 => x"80dbb404",
  2984 => x"74902975",
  2985 => x"31701080",
  2986 => x"ee98058c",
  2987 => x"77315751",
  2988 => x"54807481",
  2989 => x"b72d9e14",
  2990 => x"ff165654",
  2991 => x"74f33802",
  2992 => x"a4050d04",
  2993 => x"02fc050d",
  2994 => x"80e6e008",
  2995 => x"135180d9",
  2996 => x"e52d80e6",
  2997 => x"e408802e",
  2998 => x"8a3880e6",
  2999 => x"e4085180",
  3000 => x"cade2d80",
  3001 => x"0b80e6e0",
  3002 => x"0c80daee",
  3003 => x"2db7ba2d",
  3004 => x"0284050d",
  3005 => x"0402fc05",
  3006 => x"0d725170",
  3007 => x"fd2eb238",
  3008 => x"70fd248b",
  3009 => x"3870fc2e",
  3010 => x"80d03880",
  3011 => x"dee40470",
  3012 => x"fe2eb938",
  3013 => x"70ff2e09",
  3014 => x"810680c8",
  3015 => x"3880e6e0",
  3016 => x"08517080",
  3017 => x"2ebe38ff",
  3018 => x"1180e6e0",
  3019 => x"0c80dee4",
  3020 => x"0480e6e0",
  3021 => x"08f00570",
  3022 => x"80e6e00c",
  3023 => x"51708025",
  3024 => x"a338800b",
  3025 => x"80e6e00c",
  3026 => x"80dee404",
  3027 => x"80e6e008",
  3028 => x"810580e6",
  3029 => x"e00c80de",
  3030 => x"e40480e6",
  3031 => x"e0089005",
  3032 => x"80e6e00c",
  3033 => x"80daee2d",
  3034 => x"b7ba2d02",
  3035 => x"84050d04",
  3036 => x"02fc050d",
  3037 => x"800b80e6",
  3038 => x"e00c80da",
  3039 => x"ee2db6c3",
  3040 => x"2d80e6e4",
  3041 => x"0880e6d0",
  3042 => x"0c80e5ac",
  3043 => x"51b8e02d",
  3044 => x"0284050d",
  3045 => x"047180ee",
  3046 => x"940c0400",
  3047 => x"00ffffff",
  3048 => x"ff00ffff",
  3049 => x"ffff00ff",
  3050 => x"ffffff00",
  3051 => x"52657365",
  3052 => x"7420496e",
  3053 => x"74656c6c",
  3054 => x"69766973",
  3055 => x"696f6e00",
  3056 => x"53776170",
  3057 => x"206a6f79",
  3058 => x"73746963",
  3059 => x"6b730000",
  3060 => x"5363616e",
  3061 => x"6c696e65",
  3062 => x"73000000",
  3063 => x"4c6f6164",
  3064 => x"20524f4d",
  3065 => x"20100000",
  3066 => x"45786974",
  3067 => x"00000000",
  3068 => x"524f4d20",
  3069 => x"4d617020",
  3070 => x"74797065",
  3071 => x"20417574",
  3072 => x"6f000000",
  3073 => x"524f4d20",
  3074 => x"4d617020",
  3075 => x"74797065",
  3076 => x"20302020",
  3077 => x"20000000",
  3078 => x"524f4d20",
  3079 => x"4d617020",
  3080 => x"74797065",
  3081 => x"20312020",
  3082 => x"20000000",
  3083 => x"524f4d20",
  3084 => x"4d617020",
  3085 => x"74797065",
  3086 => x"20322020",
  3087 => x"20000000",
  3088 => x"524f4d20",
  3089 => x"4d617020",
  3090 => x"74797065",
  3091 => x"20332020",
  3092 => x"20000000",
  3093 => x"524f4d20",
  3094 => x"4d617020",
  3095 => x"74797065",
  3096 => x"20342020",
  3097 => x"20000000",
  3098 => x"524f4d20",
  3099 => x"4d617020",
  3100 => x"74797065",
  3101 => x"20352020",
  3102 => x"20000000",
  3103 => x"524f4d20",
  3104 => x"4d617020",
  3105 => x"74797065",
  3106 => x"20362020",
  3107 => x"20000000",
  3108 => x"524f4d20",
  3109 => x"4d617020",
  3110 => x"74797065",
  3111 => x"20372020",
  3112 => x"20000000",
  3113 => x"524f4d20",
  3114 => x"4d617020",
  3115 => x"74797065",
  3116 => x"20382020",
  3117 => x"20000000",
  3118 => x"524f4d20",
  3119 => x"4d617020",
  3120 => x"74797065",
  3121 => x"20392020",
  3122 => x"20000000",
  3123 => x"524f4d20",
  3124 => x"6c6f6164",
  3125 => x"696e6720",
  3126 => x"6661696c",
  3127 => x"65640000",
  3128 => x"4f4b0000",
  3129 => x"496e6974",
  3130 => x"69616c69",
  3131 => x"7a696e67",
  3132 => x"20534420",
  3133 => x"63617264",
  3134 => x"0a000000",
  3135 => x"16200000",
  3136 => x"14200000",
  3137 => x"15200000",
  3138 => x"53442069",
  3139 => x"6e69742e",
  3140 => x"2e2e0a00",
  3141 => x"53442063",
  3142 => x"61726420",
  3143 => x"72657365",
  3144 => x"74206661",
  3145 => x"696c6564",
  3146 => x"210a0000",
  3147 => x"53444843",
  3148 => x"20657272",
  3149 => x"6f72210a",
  3150 => x"00000000",
  3151 => x"57726974",
  3152 => x"65206661",
  3153 => x"696c6564",
  3154 => x"0a000000",
  3155 => x"52656164",
  3156 => x"20666169",
  3157 => x"6c65640a",
  3158 => x"00000000",
  3159 => x"43617264",
  3160 => x"20696e69",
  3161 => x"74206661",
  3162 => x"696c6564",
  3163 => x"0a000000",
  3164 => x"46415431",
  3165 => x"36202020",
  3166 => x"00000000",
  3167 => x"46415433",
  3168 => x"32202020",
  3169 => x"00000000",
  3170 => x"4e6f2070",
  3171 => x"61727469",
  3172 => x"74696f6e",
  3173 => x"20736967",
  3174 => x"0a000000",
  3175 => x"42616420",
  3176 => x"70617274",
  3177 => x"0a000000",
  3178 => x"4261636b",
  3179 => x"00000000",
  3180 => x"00000002",
  3181 => x"00000002",
  3182 => x"00002fac",
  3183 => x"0000035a",
  3184 => x"00000003",
  3185 => x"00003208",
  3186 => x"0000000b",
  3187 => x"00000001",
  3188 => x"00002fc0",
  3189 => x"00000002",
  3190 => x"00000001",
  3191 => x"00002fd0",
  3192 => x"00000003",
  3193 => x"00000002",
  3194 => x"00002fdc",
  3195 => x"00002f70",
  3196 => x"00000002",
  3197 => x"00002fe8",
  3198 => x"00001b60",
  3199 => x"00000000",
  3200 => x"00000000",
  3201 => x"00000000",
  3202 => x"00002ff0",
  3203 => x"00003004",
  3204 => x"00003018",
  3205 => x"0000302c",
  3206 => x"00003040",
  3207 => x"00003054",
  3208 => x"00003068",
  3209 => x"0000307c",
  3210 => x"00003090",
  3211 => x"000030a4",
  3212 => x"000030b8",
  3213 => x"00000004",
  3214 => x"000030cc",
  3215 => x"00003234",
  3216 => x"00000004",
  3217 => x"000030e0",
  3218 => x"000031b4",
  3219 => x"00000000",
  3220 => x"00000000",
  3221 => x"00000000",
  3222 => x"00000000",
  3223 => x"00000000",
  3224 => x"00000000",
  3225 => x"00000000",
  3226 => x"00000000",
  3227 => x"00000000",
  3228 => x"00000000",
  3229 => x"00000000",
  3230 => x"00000000",
  3231 => x"00000000",
  3232 => x"00000000",
  3233 => x"00000000",
  3234 => x"00000000",
  3235 => x"00000000",
  3236 => x"00000000",
  3237 => x"00000000",
  3238 => x"00000000",
  3239 => x"00000000",
  3240 => x"00000000",
  3241 => x"00000000",
  3242 => x"00000000",
  3243 => x"00000002",
  3244 => x"00003718",
  3245 => x"00002d34",
  3246 => x"00000002",
  3247 => x"00003736",
  3248 => x"00002d34",
  3249 => x"00000002",
  3250 => x"00003754",
  3251 => x"00002d34",
  3252 => x"00000002",
  3253 => x"00003772",
  3254 => x"00002d34",
  3255 => x"00000002",
  3256 => x"00003790",
  3257 => x"00002d34",
  3258 => x"00000002",
  3259 => x"000037ae",
  3260 => x"00002d34",
  3261 => x"00000002",
  3262 => x"000037cc",
  3263 => x"00002d34",
  3264 => x"00000002",
  3265 => x"000037ea",
  3266 => x"00002d34",
  3267 => x"00000002",
  3268 => x"00003808",
  3269 => x"00002d34",
  3270 => x"00000002",
  3271 => x"00003826",
  3272 => x"00002d34",
  3273 => x"00000002",
  3274 => x"00003844",
  3275 => x"00002d34",
  3276 => x"00000002",
  3277 => x"00003862",
  3278 => x"00002d34",
  3279 => x"00000002",
  3280 => x"00003880",
  3281 => x"00002d34",
  3282 => x"00000004",
  3283 => x"000031a8",
  3284 => x"00000000",
  3285 => x"00000000",
  3286 => x"00000000",
  3287 => x"00002ef5",
  3288 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

