library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity ASTEROIDS_PROG_ROM_0 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of ASTEROIDS_PROG_ROM_0 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"4C",X"F3",X"7C",X"20",X"FA",X"6E",X"20",X"D8",X"6E",X"20",X"68",X"71",X"AD",X"07",X"20",X"30",
		X"FE",X"46",X"5B",X"90",X"F7",X"AD",X"02",X"20",X"30",X"FB",X"AD",X"01",X"40",X"49",X"02",X"8D",
		X"01",X"40",X"8D",X"00",X"30",X"8D",X"00",X"34",X"E6",X"5C",X"D0",X"02",X"E6",X"5D",X"A2",X"40",
		X"29",X"02",X"D0",X"02",X"A2",X"44",X"A9",X"02",X"85",X"02",X"86",X"03",X"20",X"85",X"68",X"B0",
		X"C2",X"20",X"5C",X"76",X"20",X"90",X"6D",X"10",X"1B",X"20",X"C4",X"73",X"B0",X"16",X"A5",X"5A",
		X"D0",X"0C",X"20",X"D7",X"6C",X"20",X"74",X"6E",X"20",X"3F",X"70",X"20",X"93",X"6B",X"20",X"57",
		X"6F",X"20",X"F0",X"69",X"20",X"4F",X"72",X"20",X"55",X"75",X"A9",X"7F",X"AA",X"20",X"03",X"7C",
		X"20",X"B5",X"77",X"20",X"C0",X"7B",X"AD",X"FB",X"02",X"F0",X"03",X"CE",X"FB",X"02",X"0D",X"F6",
		X"02",X"D0",X"89",X"F0",X"84",X"A5",X"1C",X"F0",X"14",X"A5",X"5A",X"D0",X"03",X"4C",X"60",X"69",
		X"C6",X"5A",X"20",X"E2",X"69",X"18",X"60",X"A9",X"02",X"85",X"70",X"D0",X"13",X"A5",X"71",X"29",
		X"03",X"F0",X"F4",X"18",X"69",X"07",X"A8",X"A5",X"32",X"25",X"33",X"10",X"03",X"20",X"F6",X"77",
		X"A4",X"70",X"F0",X"E1",X"A2",X"01",X"AD",X"03",X"24",X"30",X"23",X"C0",X"02",X"90",X"7C",X"AD",
		X"04",X"24",X"10",X"77",X"A5",X"6F",X"09",X"04",X"85",X"6F",X"8D",X"00",X"32",X"20",X"D8",X"6E",
		X"20",X"68",X"71",X"20",X"E8",X"71",X"A5",X"56",X"85",X"58",X"A2",X"02",X"C6",X"70",X"86",X"1C",
		X"C6",X"70",X"A5",X"6F",X"29",X"F8",X"45",X"1C",X"85",X"6F",X"8D",X"00",X"32",X"20",X"E8",X"71",
		X"A9",X"01",X"8D",X"FA",X"02",X"8D",X"FA",X"03",X"A9",X"92",X"8D",X"F8",X"02",X"8D",X"F8",X"03",
		X"8D",X"F7",X"03",X"8D",X"F7",X"02",X"A9",X"7F",X"8D",X"FB",X"02",X"8D",X"FB",X"03",X"A9",X"05",
		X"8D",X"FD",X"02",X"8D",X"FD",X"03",X"A9",X"FF",X"85",X"32",X"85",X"33",X"A9",X"80",X"85",X"5A",
		X"0A",X"85",X"18",X"85",X"19",X"A5",X"56",X"85",X"57",X"A9",X"04",X"85",X"6C",X"85",X"6E",X"A9",
		X"30",X"8D",X"FC",X"02",X"8D",X"FC",X"03",X"8D",X"00",X"3E",X"60",X"A5",X"32",X"25",X"32",X"10",
		X"0B",X"A5",X"5C",X"29",X"20",X"D0",X"05",X"A0",X"06",X"20",X"F6",X"77",X"A5",X"5C",X"29",X"0F",
		X"D0",X"0C",X"A9",X"01",X"C5",X"70",X"69",X"01",X"49",X"01",X"45",X"6F",X"85",X"6F",X"18",X"60",
		X"A5",X"5C",X"29",X"3F",X"D0",X"0A",X"AD",X"FC",X"02",X"C9",X"08",X"F0",X"03",X"CE",X"FC",X"02",
		X"A6",X"18",X"B5",X"57",X"D0",X"1C",X"AD",X"1F",X"02",X"0D",X"20",X"02",X"0D",X"21",X"02",X"0D",
		X"22",X"02",X"D0",X"0E",X"A0",X"07",X"20",X"F6",X"77",X"A5",X"1C",X"C9",X"02",X"90",X"03",X"20",
		X"E2",X"69",X"AD",X"1B",X"02",X"D0",X"36",X"AD",X"FA",X"02",X"C9",X"80",X"D0",X"2F",X"A9",X"10",
		X"8D",X"FA",X"02",X"A6",X"1C",X"A5",X"57",X"05",X"58",X"F0",X"24",X"20",X"2D",X"70",X"CA",X"F0",
		X"1C",X"A9",X"80",X"85",X"5A",X"A5",X"18",X"49",X"01",X"AA",X"B5",X"57",X"F0",X"0F",X"86",X"18",
		X"A9",X"04",X"45",X"6F",X"85",X"6F",X"8D",X"00",X"32",X"8A",X"0A",X"85",X"19",X"18",X"60",X"86",
		X"1A",X"A9",X"FF",X"85",X"1C",X"20",X"FA",X"6E",X"A5",X"6F",X"29",X"F8",X"09",X"03",X"85",X"6F",
		X"18",X"60",X"A0",X"01",X"20",X"F6",X"77",X"A4",X"18",X"C8",X"98",X"20",X"D1",X"7B",X"60",X"62",
		X"A2",X"07",X"BD",X"1B",X"02",X"F0",X"02",X"10",X"04",X"CA",X"10",X"F6",X"60",X"A0",X"1C",X"E0",
		X"04",X"B0",X"07",X"88",X"8A",X"D0",X"03",X"88",X"30",X"EF",X"B9",X"00",X"02",X"F0",X"F8",X"30",
		X"F6",X"85",X"0B",X"B9",X"AF",X"02",X"38",X"FD",X"CA",X"02",X"85",X"08",X"B9",X"69",X"02",X"FD",
		X"84",X"02",X"4A",X"66",X"08",X"0A",X"F0",X"0C",X"10",X"6D",X"49",X"FE",X"D0",X"69",X"A5",X"08",
		X"49",X"FF",X"85",X"08",X"B9",X"D2",X"02",X"38",X"FD",X"ED",X"02",X"85",X"09",X"B9",X"8C",X"02",
		X"FD",X"A7",X"02",X"4A",X"66",X"09",X"0A",X"F0",X"0C",X"10",X"4C",X"49",X"FE",X"D0",X"48",X"A5",
		X"09",X"49",X"FF",X"85",X"09",X"A9",X"2A",X"46",X"0B",X"B0",X"08",X"A9",X"48",X"46",X"0B",X"B0",
		X"02",X"A9",X"84",X"E0",X"01",X"B0",X"02",X"69",X"1C",X"D0",X"0C",X"69",X"12",X"AE",X"1C",X"02",
		X"CA",X"F0",X"02",X"69",X"12",X"A2",X"01",X"C5",X"08",X"90",X"1C",X"C5",X"09",X"90",X"18",X"85",
		X"0B",X"4A",X"18",X"65",X"0B",X"85",X"0B",X"A5",X"09",X"65",X"08",X"B0",X"0A",X"C5",X"0B",X"B0",
		X"06",X"20",X"0F",X"6B",X"4C",X"F9",X"69",X"88",X"30",X"FA",X"4C",X"0A",X"6A",X"B9",X"00",X"02",
		X"29",X"07",X"85",X"08",X"20",X"B5",X"77",X"29",X"18",X"05",X"08",X"9D",X"00",X"02",X"B9",X"AF",
		X"02",X"9D",X"AF",X"02",X"B9",X"69",X"02",X"9D",X"69",X"02",X"B9",X"D2",X"02",X"9D",X"D2",X"02",
		X"B9",X"8C",X"02",X"9D",X"8C",X"02",X"B9",X"23",X"02",X"9D",X"23",X"02",X"B9",X"46",X"02",X"9D",
		X"46",X"02",X"60",X"85",X"0B",X"86",X"0C",X"A0",X"00",X"C8",X"B1",X"0B",X"45",X"09",X"91",X"02",
		X"88",X"C9",X"F0",X"B0",X"1E",X"C9",X"A0",X"B0",X"16",X"B1",X"0B",X"91",X"02",X"C8",X"C8",X"B1",
		X"0B",X"91",X"02",X"C8",X"B1",X"0B",X"45",X"08",X"65",X"17",X"91",X"02",X"C8",X"D0",X"DA",X"88",
		X"4C",X"39",X"7C",X"B1",X"0B",X"45",X"08",X"18",X"65",X"17",X"91",X"02",X"C8",X"D0",X"ED",X"E0",
		X"01",X"D0",X"08",X"C0",X"1B",X"D0",X"12",X"A2",X"00",X"A0",X"1C",X"8A",X"D0",X"1E",X"A9",X"81",
		X"8D",X"FA",X"02",X"A6",X"18",X"D6",X"57",X"A2",X"00",X"A9",X"A0",X"9D",X"1B",X"02",X"A9",X"00",
		X"9D",X"3E",X"02",X"9D",X"61",X"02",X"C0",X"1B",X"90",X"0D",X"B0",X"37",X"A9",X"00",X"9D",X"1B",
		X"02",X"C0",X"1B",X"F0",X"21",X"B0",X"2C",X"20",X"EC",X"75",X"B9",X"00",X"02",X"29",X"03",X"49",
		X"02",X"4A",X"6A",X"6A",X"09",X"3F",X"85",X"69",X"A9",X"A0",X"99",X"00",X"02",X"A9",X"00",X"99",
		X"23",X"02",X"99",X"46",X"02",X"60",X"8A",X"A6",X"18",X"D6",X"57",X"AA",X"A9",X"81",X"8D",X"FA",
		X"02",X"D0",X"D7",X"AD",X"F8",X"02",X"8D",X"F7",X"02",X"A5",X"1C",X"F0",X"CD",X"86",X"0D",X"A6",
		X"19",X"AD",X"1C",X"02",X"4A",X"A9",X"99",X"B0",X"02",X"A9",X"20",X"20",X"97",X"73",X"A6",X"0D",
		X"4C",X"4A",X"6B",X"A5",X"5C",X"29",X"03",X"F0",X"01",X"60",X"AD",X"1C",X"02",X"30",X"FA",X"F0",
		X"03",X"4C",X"34",X"6C",X"A5",X"1C",X"F0",X"07",X"AD",X"1B",X"02",X"F0",X"EC",X"30",X"EA",X"AD",
		X"F9",X"02",X"F0",X"03",X"CE",X"F9",X"02",X"CE",X"F7",X"02",X"D0",X"DD",X"A9",X"01",X"8D",X"F7",
		X"02",X"AD",X"F9",X"02",X"F0",X"0A",X"AD",X"F6",X"02",X"F0",X"CE",X"CD",X"FD",X"02",X"B0",X"C9",
		X"AD",X"F8",X"02",X"38",X"E9",X"06",X"C9",X"20",X"90",X"03",X"8D",X"F8",X"02",X"A9",X"00",X"8D",
		X"CB",X"02",X"8D",X"85",X"02",X"20",X"B5",X"77",X"4A",X"6E",X"EE",X"02",X"4A",X"6E",X"EE",X"02",
		X"4A",X"6E",X"EE",X"02",X"C9",X"18",X"90",X"02",X"29",X"17",X"8D",X"A8",X"02",X"A2",X"10",X"24",
		X"60",X"70",X"0C",X"A9",X"1F",X"8D",X"85",X"02",X"A9",X"FF",X"8D",X"CB",X"02",X"A2",X"F0",X"8E",
		X"3F",X"02",X"A2",X"02",X"AD",X"F8",X"02",X"30",X"17",X"A4",X"19",X"B9",X"53",X"00",X"C9",X"30",
		X"B0",X"0D",X"20",X"B5",X"77",X"85",X"08",X"AD",X"F8",X"02",X"4A",X"C5",X"08",X"B0",X"01",X"CA",
		X"8E",X"1C",X"02",X"60",X"A5",X"5C",X"0A",X"D0",X"0C",X"20",X"B5",X"77",X"29",X"03",X"AA",X"BD",
		X"D1",X"6C",X"8D",X"62",X"02",X"A5",X"1C",X"F0",X"05",X"AD",X"FA",X"02",X"D0",X"05",X"CE",X"F7",
		X"02",X"F0",X"01",X"60",X"A9",X"0A",X"8D",X"F7",X"02",X"AD",X"1C",X"02",X"4A",X"F0",X"06",X"20",
		X"B5",X"77",X"4C",X"C2",X"6C",X"AD",X"3F",X"02",X"C9",X"80",X"6A",X"85",X"0C",X"AD",X"CA",X"02",
		X"38",X"ED",X"CB",X"02",X"85",X"0B",X"AD",X"84",X"02",X"ED",X"85",X"02",X"20",X"EC",X"77",X"C9",
		X"40",X"90",X"06",X"C9",X"C0",X"B0",X"02",X"49",X"FF",X"AA",X"AD",X"62",X"02",X"C9",X"80",X"6A",
		X"85",X"0C",X"AD",X"ED",X"02",X"38",X"ED",X"EE",X"02",X"85",X"0B",X"AD",X"A7",X"02",X"ED",X"A8",
		X"02",X"20",X"EC",X"77",X"A8",X"20",X"F0",X"76",X"85",X"62",X"20",X"B5",X"77",X"A6",X"19",X"B4",
		X"53",X"C0",X"35",X"A2",X"00",X"90",X"01",X"E8",X"3D",X"CD",X"6C",X"10",X"03",X"1D",X"CF",X"6C",
		X"65",X"62",X"85",X"62",X"A0",X"03",X"A2",X"01",X"86",X"0E",X"4C",X"F2",X"6C",X"8F",X"87",X"70",
		X"78",X"F0",X"00",X"00",X"10",X"00",X"00",X"A5",X"1C",X"F0",X"21",X"0E",X"04",X"20",X"66",X"63",
		X"24",X"63",X"10",X"18",X"70",X"16",X"AD",X"FA",X"02",X"D0",X"11",X"AA",X"A9",X"03",X"85",X"0E",
		X"A0",X"07",X"B9",X"1B",X"02",X"F0",X"06",X"88",X"C4",X"0E",X"D0",X"F6",X"60",X"86",X"0D",X"A9",
		X"12",X"99",X"1B",X"02",X"B5",X"61",X"20",X"D2",X"77",X"A6",X"0D",X"C9",X"80",X"6A",X"85",X"09",
		X"18",X"7D",X"3E",X"02",X"30",X"08",X"C9",X"70",X"90",X"0A",X"A9",X"6F",X"D0",X"06",X"C9",X"91",
		X"B0",X"02",X"A9",X"91",X"99",X"3E",X"02",X"B5",X"61",X"20",X"D5",X"77",X"A6",X"0D",X"C9",X"80",
		X"6A",X"85",X"0C",X"18",X"7D",X"61",X"02",X"30",X"08",X"C9",X"70",X"90",X"0A",X"A9",X"6F",X"D0",
		X"06",X"C9",X"91",X"B0",X"02",X"A9",X"91",X"99",X"61",X"02",X"A2",X"00",X"A5",X"09",X"10",X"01",
		X"CA",X"86",X"08",X"A6",X"0D",X"C9",X"80",X"6A",X"18",X"65",X"09",X"18",X"7D",X"CA",X"02",X"99",
		X"CA",X"02",X"A5",X"08",X"7D",X"84",X"02",X"99",X"84",X"02",X"A2",X"00",X"A5",X"0C",X"10",X"01",
		X"CA",X"86",X"0B",X"A6",X"0D",X"C9",X"80",X"6A",X"18",X"65",X"0C",X"18",X"7D",X"ED",X"02",X"99",
		X"ED",X"02",X"A5",X"0B",X"7D",X"A7",X"02",X"99",X"A7",X"02",X"A9",X"80",X"95",X"66",X"60",X"D6",
		X"A5",X"32",X"25",X"33",X"10",X"01",X"60",X"A5",X"1A",X"4A",X"F0",X"18",X"A0",X"01",X"20",X"F6",
		X"77",X"A0",X"02",X"A6",X"33",X"10",X"01",X"88",X"84",X"18",X"A5",X"5C",X"29",X"10",X"D0",X"04",
		X"98",X"20",X"D1",X"7B",X"46",X"18",X"20",X"B2",X"73",X"A0",X"02",X"20",X"F6",X"77",X"A0",X"03",
		X"20",X"F6",X"77",X"A0",X"04",X"20",X"F6",X"77",X"A0",X"05",X"20",X"F6",X"77",X"A9",X"20",X"85",
		X"00",X"A9",X"64",X"A2",X"39",X"20",X"03",X"7C",X"A9",X"70",X"20",X"DE",X"7C",X"A6",X"18",X"B4",
		X"32",X"84",X"0B",X"98",X"18",X"65",X"31",X"85",X"0C",X"20",X"1A",X"6F",X"A4",X"0B",X"C8",X"20",
		X"1A",X"6F",X"A4",X"0B",X"C8",X"C8",X"20",X"1A",X"6F",X"AD",X"03",X"20",X"2A",X"26",X"63",X"A5",
		X"63",X"29",X"1F",X"C9",X"07",X"D0",X"27",X"E6",X"31",X"A5",X"31",X"C9",X"03",X"90",X"13",X"A6",
		X"18",X"A9",X"FF",X"95",X"32",X"A2",X"00",X"86",X"18",X"86",X"31",X"A2",X"F0",X"86",X"5D",X"4C",
		X"B2",X"73",X"E6",X"0C",X"A6",X"0C",X"A9",X"F4",X"85",X"5D",X"A9",X"0B",X"95",X"34",X"A5",X"5D",
		X"D0",X"08",X"A9",X"FF",X"85",X"32",X"85",X"33",X"30",X"DB",X"A5",X"5C",X"29",X"07",X"D0",X"31",
		X"AD",X"07",X"24",X"10",X"04",X"A9",X"01",X"D0",X"07",X"AD",X"06",X"24",X"10",X"23",X"A9",X"FF",
		X"A6",X"0C",X"18",X"75",X"34",X"30",X"10",X"C9",X"0B",X"B0",X"0E",X"C9",X"01",X"F0",X"04",X"A9",
		X"00",X"F0",X"0C",X"A9",X"0B",X"D0",X"08",X"A9",X"24",X"C9",X"25",X"90",X"02",X"A9",X"00",X"95",
		X"34",X"A9",X"00",X"60",X"A5",X"1C",X"F0",X"5F",X"AD",X"1B",X"02",X"30",X"5A",X"AD",X"FA",X"02",
		X"D0",X"55",X"AD",X"03",X"20",X"10",X"50",X"A9",X"00",X"8D",X"1B",X"02",X"8D",X"3E",X"02",X"8D",
		X"61",X"02",X"A9",X"30",X"8D",X"FA",X"02",X"20",X"B5",X"77",X"29",X"1F",X"C9",X"1D",X"90",X"02",
		X"A9",X"1C",X"C9",X"03",X"B0",X"02",X"A9",X"03",X"8D",X"84",X"02",X"A2",X"05",X"20",X"B5",X"77",
		X"CA",X"D0",X"FA",X"29",X"1F",X"E8",X"C9",X"18",X"90",X"0C",X"29",X"07",X"0A",X"69",X"04",X"CD",
		X"F6",X"02",X"90",X"02",X"A2",X"80",X"C9",X"15",X"90",X"02",X"A9",X"14",X"C9",X"03",X"B0",X"02",
		X"A9",X"03",X"8D",X"A7",X"02",X"86",X"59",X"60",X"A9",X"02",X"8D",X"F5",X"02",X"A2",X"03",X"4E",
		X"02",X"28",X"B0",X"01",X"E8",X"86",X"56",X"A9",X"00",X"A2",X"03",X"9D",X"1B",X"02",X"9D",X"1F",
		X"02",X"95",X"52",X"CA",X"10",X"F5",X"8D",X"F6",X"02",X"60",X"A9",X"00",X"8D",X"00",X"36",X"8D",
		X"00",X"3A",X"8D",X"00",X"3C",X"8D",X"01",X"3C",X"8D",X"03",X"3C",X"8D",X"04",X"3C",X"8D",X"05",
		X"3C",X"85",X"69",X"85",X"66",X"85",X"67",X"85",X"68",X"60",X"B9",X"34",X"00",X"0A",X"A8",X"D0",
		X"14",X"A5",X"32",X"25",X"33",X"30",X"0E",X"A9",X"72",X"A2",X"F8",X"20",X"45",X"7D",X"A9",X"01",
		X"A2",X"F8",X"4C",X"45",X"7D",X"BE",X"D5",X"56",X"B9",X"D4",X"56",X"4C",X"45",X"7D",X"F0",X"16",
		X"84",X"08",X"A2",X"D5",X"A0",X"E0",X"84",X"00",X"20",X"03",X"7C",X"A2",X"DA",X"A9",X"54",X"20",
		X"FC",X"7B",X"C6",X"08",X"D0",X"F5",X"60",X"A2",X"22",X"BD",X"00",X"02",X"D0",X"04",X"CA",X"10",
		X"F8",X"60",X"10",X"63",X"20",X"08",X"77",X"4A",X"4A",X"4A",X"4A",X"E0",X"1B",X"D0",X"07",X"A5",
		X"5C",X"29",X"01",X"4A",X"F0",X"01",X"38",X"7D",X"00",X"02",X"30",X"25",X"E0",X"1B",X"F0",X"13",
		X"B0",X"17",X"CE",X"F6",X"02",X"D0",X"05",X"A0",X"7F",X"8C",X"FB",X"02",X"A9",X"00",X"9D",X"00",
		X"02",X"F0",X"CB",X"20",X"E8",X"71",X"4C",X"8C",X"6F",X"AD",X"F8",X"02",X"8D",X"F7",X"02",X"D0",
		X"EB",X"9D",X"00",X"02",X"29",X"F0",X"18",X"69",X"10",X"E0",X"1B",X"D0",X"02",X"A9",X"00",X"A8",
		X"BD",X"AF",X"02",X"85",X"04",X"BD",X"69",X"02",X"85",X"05",X"BD",X"D2",X"02",X"85",X"06",X"BD",
		X"8C",X"02",X"85",X"07",X"4C",X"27",X"70",X"18",X"A0",X"00",X"BD",X"23",X"02",X"10",X"01",X"88",
		X"7D",X"AF",X"02",X"9D",X"AF",X"02",X"85",X"04",X"98",X"7D",X"69",X"02",X"C9",X"20",X"90",X"0C",
		X"29",X"1F",X"E0",X"1C",X"D0",X"06",X"20",X"2D",X"70",X"4C",X"5E",X"6F",X"9D",X"69",X"02",X"85",
		X"05",X"18",X"A0",X"00",X"BD",X"46",X"02",X"10",X"02",X"A0",X"FF",X"7D",X"D2",X"02",X"9D",X"D2");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
