-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80e6",
     9 => x"8c080b0b",
    10 => x"80e69008",
    11 => x"0b0b80e6",
    12 => x"94080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"e6940c0b",
    16 => x"0b80e690",
    17 => x"0c0b0b80",
    18 => x"e68c0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80dfc8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80e68c70",
    57 => x"80f0c827",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c51b192",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80e6",
    65 => x"9c0c9f0b",
    66 => x"80e6a00c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"e6a008ff",
    70 => x"0580e6a0",
    71 => x"0c80e6a0",
    72 => x"088025e8",
    73 => x"3880e69c",
    74 => x"08ff0580",
    75 => x"e69c0c80",
    76 => x"e69c0880",
    77 => x"25d03880",
    78 => x"0b80e6a0",
    79 => x"0c800b80",
    80 => x"e69c0c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80e69c08",
   100 => x"25913882",
   101 => x"c82d80e6",
   102 => x"9c08ff05",
   103 => x"80e69c0c",
   104 => x"838a0480",
   105 => x"e69c0880",
   106 => x"e6a00853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80e69c08",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"e6a00881",
   116 => x"0580e6a0",
   117 => x"0c80e6a0",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80e6a0",
   121 => x"0c80e69c",
   122 => x"08810580",
   123 => x"e69c0c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480e6",
   128 => x"a0088105",
   129 => x"80e6a00c",
   130 => x"80e6a008",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80e6a0",
   134 => x"0c80e69c",
   135 => x"08810580",
   136 => x"e69c0c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"e6a40cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565481ff",
   169 => x"06527372",
   170 => x"25893871",
   171 => x"54820b80",
   172 => x"e6a40c72",
   173 => x"882c7381",
   174 => x"ff065455",
   175 => x"7473258d",
   176 => x"387280e6",
   177 => x"a4088407",
   178 => x"80e6a40c",
   179 => x"5573842b",
   180 => x"86a07125",
   181 => x"83713170",
   182 => x"0b0b80e2",
   183 => x"e00c8171",
   184 => x"2bff05f6",
   185 => x"880cfdfc",
   186 => x"13ff122c",
   187 => x"788829ff",
   188 => x"94057081",
   189 => x"2c80e6a4",
   190 => x"08525852",
   191 => x"55515254",
   192 => x"76802e85",
   193 => x"38708107",
   194 => x"5170f694",
   195 => x"0c710981",
   196 => x"05f6800c",
   197 => x"72098105",
   198 => x"f6840c02",
   199 => x"94050d04",
   200 => x"02f4050d",
   201 => x"74537270",
   202 => x"81055480",
   203 => x"f52d5271",
   204 => x"802e8938",
   205 => x"71518384",
   206 => x"2d86a604",
   207 => x"810b80e6",
   208 => x"8c0c028c",
   209 => x"050d0402",
   210 => x"fc050d81",
   211 => x"808051c0",
   212 => x"115170fb",
   213 => x"38028405",
   214 => x"0d0402fc",
   215 => x"050dec51",
   216 => x"83710c86",
   217 => x"c72d8271",
   218 => x"0c028405",
   219 => x"0d0402fc",
   220 => x"050dec51",
   221 => x"8a710c86",
   222 => x"c72d86c7",
   223 => x"2d86c72d",
   224 => x"86c72d86",
   225 => x"c72d86c7",
   226 => x"2d86c72d",
   227 => x"86c72d86",
   228 => x"c72d86c7",
   229 => x"2d86c72d",
   230 => x"86c72d86",
   231 => x"c72d86c7",
   232 => x"2d86c72d",
   233 => x"86c72d86",
   234 => x"c72d86c7",
   235 => x"2d86c72d",
   236 => x"86c72d86",
   237 => x"c72d86c7",
   238 => x"2d86c72d",
   239 => x"86c72d86",
   240 => x"c72d86c7",
   241 => x"2d86c72d",
   242 => x"86c72d86",
   243 => x"c72d86c7",
   244 => x"2d86c72d",
   245 => x"86c72d86",
   246 => x"c72d86c7",
   247 => x"2d86c72d",
   248 => x"86c72d86",
   249 => x"c72d86c7",
   250 => x"2d86c72d",
   251 => x"86c72d86",
   252 => x"c72d86c7",
   253 => x"2d86c72d",
   254 => x"86c72d86",
   255 => x"c72d86c7",
   256 => x"2d86c72d",
   257 => x"86c72d86",
   258 => x"c72d86c7",
   259 => x"2d86c72d",
   260 => x"86c72d86",
   261 => x"c72d86c7",
   262 => x"2d86c72d",
   263 => x"86c72d86",
   264 => x"c72d86c7",
   265 => x"2d86c72d",
   266 => x"86c72d86",
   267 => x"c72d86c7",
   268 => x"2d86c72d",
   269 => x"86c72d86",
   270 => x"c72d86c7",
   271 => x"2d86c72d",
   272 => x"86c72d86",
   273 => x"c72d86c7",
   274 => x"2d86c72d",
   275 => x"86c72d86",
   276 => x"c72d86c7",
   277 => x"2d86c72d",
   278 => x"86c72d86",
   279 => x"c72d86c7",
   280 => x"2d86c72d",
   281 => x"86c72d86",
   282 => x"c72d86c7",
   283 => x"2d86c72d",
   284 => x"86c72d86",
   285 => x"c72d86c7",
   286 => x"2d86c72d",
   287 => x"86c72d86",
   288 => x"c72d86c7",
   289 => x"2d86c72d",
   290 => x"86c72d86",
   291 => x"c72d86c7",
   292 => x"2d86c72d",
   293 => x"86c72d86",
   294 => x"c72d86c7",
   295 => x"2d86c72d",
   296 => x"86c72d86",
   297 => x"c72d86c7",
   298 => x"2d86c72d",
   299 => x"86c72d86",
   300 => x"c72d86c7",
   301 => x"2d86c72d",
   302 => x"86c72d86",
   303 => x"c72d86c7",
   304 => x"2d86c72d",
   305 => x"86c72d86",
   306 => x"c72d86c7",
   307 => x"2d86c72d",
   308 => x"86c72d86",
   309 => x"c72d86c7",
   310 => x"2d86c72d",
   311 => x"86c72d86",
   312 => x"c72d86c7",
   313 => x"2d86c72d",
   314 => x"86c72d86",
   315 => x"c72d86c7",
   316 => x"2d86c72d",
   317 => x"86c72d86",
   318 => x"c72d86c7",
   319 => x"2d86c72d",
   320 => x"86c72d86",
   321 => x"c72d86c7",
   322 => x"2d86c72d",
   323 => x"86c72d86",
   324 => x"c72d86c7",
   325 => x"2d86c72d",
   326 => x"86c72d86",
   327 => x"c72d86c7",
   328 => x"2d86c72d",
   329 => x"86c72d86",
   330 => x"c72d86c7",
   331 => x"2d86c72d",
   332 => x"86c72d86",
   333 => x"c72d86c7",
   334 => x"2d86c72d",
   335 => x"86c72d86",
   336 => x"c72d86c7",
   337 => x"2d86c72d",
   338 => x"86c72d86",
   339 => x"c72d86c7",
   340 => x"2d86c72d",
   341 => x"86c72d86",
   342 => x"c72d86c7",
   343 => x"2d86c72d",
   344 => x"86c72d86",
   345 => x"c72d86c7",
   346 => x"2d86c72d",
   347 => x"86c72d86",
   348 => x"c72d86c7",
   349 => x"2d86c72d",
   350 => x"86c72d86",
   351 => x"c72d86c7",
   352 => x"2d86c72d",
   353 => x"86c72d86",
   354 => x"c72d86c7",
   355 => x"2d86c72d",
   356 => x"86c72d86",
   357 => x"c72d86c7",
   358 => x"2d86c72d",
   359 => x"86c72d86",
   360 => x"c72d86c7",
   361 => x"2d86c72d",
   362 => x"86c72d86",
   363 => x"c72d86c7",
   364 => x"2d86c72d",
   365 => x"86c72d86",
   366 => x"c72d86c7",
   367 => x"2d86c72d",
   368 => x"86c72d86",
   369 => x"c72d86c7",
   370 => x"2d86c72d",
   371 => x"86c72d86",
   372 => x"c72d86c7",
   373 => x"2d86c72d",
   374 => x"86c72d86",
   375 => x"c72d86c7",
   376 => x"2d86c72d",
   377 => x"86c72d86",
   378 => x"c72d86c7",
   379 => x"2d86c72d",
   380 => x"86c72d86",
   381 => x"c72d86c7",
   382 => x"2d86c72d",
   383 => x"86c72d86",
   384 => x"c72d86c7",
   385 => x"2d86c72d",
   386 => x"86c72d86",
   387 => x"c72d86c7",
   388 => x"2d86c72d",
   389 => x"86c72d86",
   390 => x"c72d86c7",
   391 => x"2d86c72d",
   392 => x"86c72d86",
   393 => x"c72d86c7",
   394 => x"2d86c72d",
   395 => x"86c72d86",
   396 => x"c72d86c7",
   397 => x"2d86c72d",
   398 => x"86c72d86",
   399 => x"c72d86c7",
   400 => x"2d86c72d",
   401 => x"86c72d86",
   402 => x"c72d86c7",
   403 => x"2d86c72d",
   404 => x"86c72d86",
   405 => x"c72d86c7",
   406 => x"2d86c72d",
   407 => x"86c72d86",
   408 => x"c72d86c7",
   409 => x"2d86c72d",
   410 => x"86c72d86",
   411 => x"c72d86c7",
   412 => x"2d86c72d",
   413 => x"86c72d86",
   414 => x"c72d86c7",
   415 => x"2d86c72d",
   416 => x"86c72d86",
   417 => x"c72d86c7",
   418 => x"2d86c72d",
   419 => x"86c72d86",
   420 => x"c72d86c7",
   421 => x"2d86c72d",
   422 => x"86c72d86",
   423 => x"c72d86c7",
   424 => x"2d86c72d",
   425 => x"86c72d86",
   426 => x"c72d86c7",
   427 => x"2d86c72d",
   428 => x"86c72d86",
   429 => x"c72d86c7",
   430 => x"2d86c72d",
   431 => x"86c72d86",
   432 => x"c72d86c7",
   433 => x"2d86c72d",
   434 => x"86c72d86",
   435 => x"c72d86c7",
   436 => x"2d86c72d",
   437 => x"86c72d86",
   438 => x"c72d86c7",
   439 => x"2d86c72d",
   440 => x"86c72d86",
   441 => x"c72d86c7",
   442 => x"2d86c72d",
   443 => x"86c72d86",
   444 => x"c72d86c7",
   445 => x"2d86c72d",
   446 => x"86c72d86",
   447 => x"c72d86c7",
   448 => x"2d86c72d",
   449 => x"86c72d86",
   450 => x"c72d86c7",
   451 => x"2d86c72d",
   452 => x"86c72d86",
   453 => x"c72d86c7",
   454 => x"2d86c72d",
   455 => x"86c72d86",
   456 => x"c72d86c7",
   457 => x"2d86c72d",
   458 => x"86c72d86",
   459 => x"c72d86c7",
   460 => x"2d86c72d",
   461 => x"86c72d86",
   462 => x"c72d86c7",
   463 => x"2d86c72d",
   464 => x"86c72d86",
   465 => x"c72d86c7",
   466 => x"2d86c72d",
   467 => x"86c72d86",
   468 => x"c72d86c7",
   469 => x"2d86c72d",
   470 => x"86c72d86",
   471 => x"c72d86c7",
   472 => x"2d86c72d",
   473 => x"86c72d86",
   474 => x"c72d86c7",
   475 => x"2d86c72d",
   476 => x"86c72d86",
   477 => x"c72d86c7",
   478 => x"2d86c72d",
   479 => x"86c72d86",
   480 => x"c72d86c7",
   481 => x"2d86c72d",
   482 => x"86c72d86",
   483 => x"c72d86c7",
   484 => x"2d86c72d",
   485 => x"86c72d86",
   486 => x"c72d86c7",
   487 => x"2d86c72d",
   488 => x"86c72d86",
   489 => x"c72d86c7",
   490 => x"2d86c72d",
   491 => x"86c72d86",
   492 => x"c72d86c7",
   493 => x"2d86c72d",
   494 => x"86c72d86",
   495 => x"c72d86c7",
   496 => x"2d86c72d",
   497 => x"86c72d86",
   498 => x"c72d86c7",
   499 => x"2d86c72d",
   500 => x"86c72d86",
   501 => x"c72d86c7",
   502 => x"2d86c72d",
   503 => x"86c72d86",
   504 => x"c72d86c7",
   505 => x"2d86c72d",
   506 => x"86c72d86",
   507 => x"c72d86c7",
   508 => x"2d86c72d",
   509 => x"86c72d86",
   510 => x"c72d86c7",
   511 => x"2d86c72d",
   512 => x"86c72d86",
   513 => x"c72d86c7",
   514 => x"2d86c72d",
   515 => x"86c72d86",
   516 => x"c72d86c7",
   517 => x"2d86c72d",
   518 => x"86c72d86",
   519 => x"c72d86c7",
   520 => x"2d86c72d",
   521 => x"86c72d86",
   522 => x"c72d86c7",
   523 => x"2d86c72d",
   524 => x"86c72d86",
   525 => x"c72d86c7",
   526 => x"2d86c72d",
   527 => x"86c72d86",
   528 => x"c72d86c7",
   529 => x"2d86c72d",
   530 => x"86c72d86",
   531 => x"c72d86c7",
   532 => x"2d86c72d",
   533 => x"86c72d86",
   534 => x"c72d86c7",
   535 => x"2d86c72d",
   536 => x"86c72d86",
   537 => x"c72d86c7",
   538 => x"2d86c72d",
   539 => x"86c72d86",
   540 => x"c72d86c7",
   541 => x"2d86c72d",
   542 => x"86c72d86",
   543 => x"c72d86c7",
   544 => x"2d86c72d",
   545 => x"86c72d86",
   546 => x"c72d86c7",
   547 => x"2d86c72d",
   548 => x"86c72d86",
   549 => x"c72d86c7",
   550 => x"2d86c72d",
   551 => x"86c72d86",
   552 => x"c72d86c7",
   553 => x"2d86c72d",
   554 => x"86c72d86",
   555 => x"c72d86c7",
   556 => x"2d86c72d",
   557 => x"86c72d86",
   558 => x"c72d86c7",
   559 => x"2d86c72d",
   560 => x"86c72d86",
   561 => x"c72d86c7",
   562 => x"2d86c72d",
   563 => x"86c72d86",
   564 => x"c72d86c7",
   565 => x"2d86c72d",
   566 => x"86c72d86",
   567 => x"c72d86c7",
   568 => x"2d86c72d",
   569 => x"86c72d86",
   570 => x"c72d86c7",
   571 => x"2d86c72d",
   572 => x"86c72d86",
   573 => x"c72d86c7",
   574 => x"2d86c72d",
   575 => x"86c72d86",
   576 => x"c72d86c7",
   577 => x"2d86c72d",
   578 => x"86c72d86",
   579 => x"c72d86c7",
   580 => x"2d86c72d",
   581 => x"86c72d86",
   582 => x"c72d86c7",
   583 => x"2d86c72d",
   584 => x"86c72d86",
   585 => x"c72d86c7",
   586 => x"2d86c72d",
   587 => x"86c72d86",
   588 => x"c72d86c7",
   589 => x"2d86c72d",
   590 => x"86c72d86",
   591 => x"c72d86c7",
   592 => x"2d86c72d",
   593 => x"86c72d86",
   594 => x"c72d86c7",
   595 => x"2d86c72d",
   596 => x"86c72d86",
   597 => x"c72d86c7",
   598 => x"2d86c72d",
   599 => x"86c72d86",
   600 => x"c72d86c7",
   601 => x"2d86c72d",
   602 => x"86c72d86",
   603 => x"c72d86c7",
   604 => x"2d86c72d",
   605 => x"86c72d86",
   606 => x"c72d86c7",
   607 => x"2d86c72d",
   608 => x"86c72d86",
   609 => x"c72d86c7",
   610 => x"2d86c72d",
   611 => x"86c72d86",
   612 => x"c72d86c7",
   613 => x"2d86c72d",
   614 => x"86c72d86",
   615 => x"c72d86c7",
   616 => x"2d86c72d",
   617 => x"86c72d86",
   618 => x"c72d86c7",
   619 => x"2d86c72d",
   620 => x"86c72d86",
   621 => x"c72d86c7",
   622 => x"2d86c72d",
   623 => x"86c72d86",
   624 => x"c72d86c7",
   625 => x"2d86c72d",
   626 => x"86c72d86",
   627 => x"c72d86c7",
   628 => x"2d86c72d",
   629 => x"86c72d86",
   630 => x"c72d86c7",
   631 => x"2d86c72d",
   632 => x"86c72d86",
   633 => x"c72d86c7",
   634 => x"2d86c72d",
   635 => x"86c72d86",
   636 => x"c72d86c7",
   637 => x"2d86c72d",
   638 => x"86c72d86",
   639 => x"c72d86c7",
   640 => x"2d86c72d",
   641 => x"86c72d86",
   642 => x"c72d86c7",
   643 => x"2d86c72d",
   644 => x"86c72d86",
   645 => x"c72d86c7",
   646 => x"2d86c72d",
   647 => x"86c72d86",
   648 => x"c72d86c7",
   649 => x"2d86c72d",
   650 => x"86c72d86",
   651 => x"c72d86c7",
   652 => x"2d86c72d",
   653 => x"86c72d82",
   654 => x"710c0284",
   655 => x"050d0402",
   656 => x"fc050dec",
   657 => x"5192710c",
   658 => x"86c72d86",
   659 => x"c72d86c7",
   660 => x"2d86c72d",
   661 => x"86c72d86",
   662 => x"c72d86c7",
   663 => x"2d86c72d",
   664 => x"86c72d86",
   665 => x"c72d86c7",
   666 => x"2d86c72d",
   667 => x"86c72d86",
   668 => x"c72d86c7",
   669 => x"2d86c72d",
   670 => x"86c72d86",
   671 => x"c72d86c7",
   672 => x"2d86c72d",
   673 => x"86c72d86",
   674 => x"c72d86c7",
   675 => x"2d86c72d",
   676 => x"86c72d86",
   677 => x"c72d86c7",
   678 => x"2d86c72d",
   679 => x"86c72d86",
   680 => x"c72d86c7",
   681 => x"2d86c72d",
   682 => x"86c72d86",
   683 => x"c72d86c7",
   684 => x"2d86c72d",
   685 => x"86c72d86",
   686 => x"c72d86c7",
   687 => x"2d86c72d",
   688 => x"86c72d86",
   689 => x"c72d86c7",
   690 => x"2d86c72d",
   691 => x"86c72d86",
   692 => x"c72d86c7",
   693 => x"2d86c72d",
   694 => x"86c72d86",
   695 => x"c72d86c7",
   696 => x"2d86c72d",
   697 => x"86c72d86",
   698 => x"c72d86c7",
   699 => x"2d86c72d",
   700 => x"86c72d86",
   701 => x"c72d86c7",
   702 => x"2d86c72d",
   703 => x"86c72d86",
   704 => x"c72d86c7",
   705 => x"2d86c72d",
   706 => x"86c72d86",
   707 => x"c72d86c7",
   708 => x"2d86c72d",
   709 => x"86c72d86",
   710 => x"c72d86c7",
   711 => x"2d86c72d",
   712 => x"86c72d86",
   713 => x"c72d86c7",
   714 => x"2d86c72d",
   715 => x"86c72d86",
   716 => x"c72d86c7",
   717 => x"2d86c72d",
   718 => x"86c72d86",
   719 => x"c72d86c7",
   720 => x"2d86c72d",
   721 => x"86c72d86",
   722 => x"c72d86c7",
   723 => x"2d86c72d",
   724 => x"86c72d86",
   725 => x"c72d86c7",
   726 => x"2d86c72d",
   727 => x"86c72d86",
   728 => x"c72d86c7",
   729 => x"2d86c72d",
   730 => x"86c72d86",
   731 => x"c72d86c7",
   732 => x"2d86c72d",
   733 => x"86c72d86",
   734 => x"c72d86c7",
   735 => x"2d86c72d",
   736 => x"86c72d86",
   737 => x"c72d86c7",
   738 => x"2d86c72d",
   739 => x"86c72d86",
   740 => x"c72d86c7",
   741 => x"2d86c72d",
   742 => x"86c72d86",
   743 => x"c72d86c7",
   744 => x"2d86c72d",
   745 => x"86c72d86",
   746 => x"c72d86c7",
   747 => x"2d86c72d",
   748 => x"86c72d86",
   749 => x"c72d86c7",
   750 => x"2d86c72d",
   751 => x"86c72d86",
   752 => x"c72d86c7",
   753 => x"2d86c72d",
   754 => x"86c72d86",
   755 => x"c72d86c7",
   756 => x"2d86c72d",
   757 => x"86c72d86",
   758 => x"c72d86c7",
   759 => x"2d86c72d",
   760 => x"86c72d86",
   761 => x"c72d86c7",
   762 => x"2d86c72d",
   763 => x"86c72d86",
   764 => x"c72d86c7",
   765 => x"2d86c72d",
   766 => x"86c72d86",
   767 => x"c72d86c7",
   768 => x"2d86c72d",
   769 => x"86c72d86",
   770 => x"c72d86c7",
   771 => x"2d86c72d",
   772 => x"86c72d86",
   773 => x"c72d86c7",
   774 => x"2d86c72d",
   775 => x"86c72d86",
   776 => x"c72d86c7",
   777 => x"2d86c72d",
   778 => x"86c72d86",
   779 => x"c72d86c7",
   780 => x"2d86c72d",
   781 => x"86c72d86",
   782 => x"c72d86c7",
   783 => x"2d86c72d",
   784 => x"86c72d86",
   785 => x"c72d86c7",
   786 => x"2d86c72d",
   787 => x"86c72d86",
   788 => x"c72d86c7",
   789 => x"2d86c72d",
   790 => x"86c72d86",
   791 => x"c72d86c7",
   792 => x"2d86c72d",
   793 => x"86c72d86",
   794 => x"c72d86c7",
   795 => x"2d86c72d",
   796 => x"86c72d86",
   797 => x"c72d86c7",
   798 => x"2d86c72d",
   799 => x"86c72d86",
   800 => x"c72d86c7",
   801 => x"2d86c72d",
   802 => x"86c72d86",
   803 => x"c72d86c7",
   804 => x"2d86c72d",
   805 => x"86c72d86",
   806 => x"c72d86c7",
   807 => x"2d86c72d",
   808 => x"86c72d86",
   809 => x"c72d86c7",
   810 => x"2d86c72d",
   811 => x"86c72d86",
   812 => x"c72d86c7",
   813 => x"2d86c72d",
   814 => x"86c72d86",
   815 => x"c72d86c7",
   816 => x"2d86c72d",
   817 => x"86c72d86",
   818 => x"c72d86c7",
   819 => x"2d86c72d",
   820 => x"86c72d86",
   821 => x"c72d86c7",
   822 => x"2d86c72d",
   823 => x"86c72d86",
   824 => x"c72d86c7",
   825 => x"2d86c72d",
   826 => x"86c72d86",
   827 => x"c72d86c7",
   828 => x"2d86c72d",
   829 => x"86c72d86",
   830 => x"c72d86c7",
   831 => x"2d86c72d",
   832 => x"86c72d86",
   833 => x"c72d86c7",
   834 => x"2d86c72d",
   835 => x"86c72d86",
   836 => x"c72d86c7",
   837 => x"2d86c72d",
   838 => x"86c72d86",
   839 => x"c72d86c7",
   840 => x"2d86c72d",
   841 => x"86c72d86",
   842 => x"c72d86c7",
   843 => x"2d86c72d",
   844 => x"86c72d86",
   845 => x"c72d86c7",
   846 => x"2d86c72d",
   847 => x"86c72d86",
   848 => x"c72d86c7",
   849 => x"2d86c72d",
   850 => x"86c72d86",
   851 => x"c72d86c7",
   852 => x"2d86c72d",
   853 => x"86c72d86",
   854 => x"c72d86c7",
   855 => x"2d86c72d",
   856 => x"86c72d86",
   857 => x"c72d86c7",
   858 => x"2d86c72d",
   859 => x"86c72d86",
   860 => x"c72d86c7",
   861 => x"2d86c72d",
   862 => x"86c72d86",
   863 => x"c72d86c7",
   864 => x"2d86c72d",
   865 => x"86c72d86",
   866 => x"c72d86c7",
   867 => x"2d86c72d",
   868 => x"86c72d86",
   869 => x"c72d86c7",
   870 => x"2d86c72d",
   871 => x"86c72d86",
   872 => x"c72d86c7",
   873 => x"2d86c72d",
   874 => x"86c72d86",
   875 => x"c72d86c7",
   876 => x"2d86c72d",
   877 => x"86c72d86",
   878 => x"c72d86c7",
   879 => x"2d86c72d",
   880 => x"86c72d86",
   881 => x"c72d86c7",
   882 => x"2d86c72d",
   883 => x"86c72d86",
   884 => x"c72d86c7",
   885 => x"2d86c72d",
   886 => x"86c72d86",
   887 => x"c72d86c7",
   888 => x"2d86c72d",
   889 => x"86c72d86",
   890 => x"c72d86c7",
   891 => x"2d86c72d",
   892 => x"86c72d86",
   893 => x"c72d86c7",
   894 => x"2d86c72d",
   895 => x"86c72d86",
   896 => x"c72d86c7",
   897 => x"2d86c72d",
   898 => x"86c72d86",
   899 => x"c72d86c7",
   900 => x"2d86c72d",
   901 => x"86c72d86",
   902 => x"c72d86c7",
   903 => x"2d86c72d",
   904 => x"86c72d86",
   905 => x"c72d86c7",
   906 => x"2d86c72d",
   907 => x"86c72d86",
   908 => x"c72d86c7",
   909 => x"2d86c72d",
   910 => x"86c72d86",
   911 => x"c72d86c7",
   912 => x"2d86c72d",
   913 => x"86c72d86",
   914 => x"c72d86c7",
   915 => x"2d86c72d",
   916 => x"86c72d86",
   917 => x"c72d86c7",
   918 => x"2d86c72d",
   919 => x"86c72d86",
   920 => x"c72d86c7",
   921 => x"2d86c72d",
   922 => x"86c72d86",
   923 => x"c72d86c7",
   924 => x"2d86c72d",
   925 => x"86c72d86",
   926 => x"c72d86c7",
   927 => x"2d86c72d",
   928 => x"86c72d86",
   929 => x"c72d86c7",
   930 => x"2d86c72d",
   931 => x"86c72d86",
   932 => x"c72d86c7",
   933 => x"2d86c72d",
   934 => x"86c72d86",
   935 => x"c72d86c7",
   936 => x"2d86c72d",
   937 => x"86c72d86",
   938 => x"c72d86c7",
   939 => x"2d86c72d",
   940 => x"86c72d86",
   941 => x"c72d86c7",
   942 => x"2d86c72d",
   943 => x"86c72d86",
   944 => x"c72d86c7",
   945 => x"2d86c72d",
   946 => x"86c72d86",
   947 => x"c72d86c7",
   948 => x"2d86c72d",
   949 => x"86c72d86",
   950 => x"c72d86c7",
   951 => x"2d86c72d",
   952 => x"86c72d86",
   953 => x"c72d86c7",
   954 => x"2d86c72d",
   955 => x"86c72d86",
   956 => x"c72d86c7",
   957 => x"2d86c72d",
   958 => x"86c72d86",
   959 => x"c72d86c7",
   960 => x"2d86c72d",
   961 => x"86c72d86",
   962 => x"c72d86c7",
   963 => x"2d86c72d",
   964 => x"86c72d86",
   965 => x"c72d86c7",
   966 => x"2d86c72d",
   967 => x"86c72d86",
   968 => x"c72d86c7",
   969 => x"2d86c72d",
   970 => x"86c72d86",
   971 => x"c72d86c7",
   972 => x"2d86c72d",
   973 => x"86c72d86",
   974 => x"c72d86c7",
   975 => x"2d86c72d",
   976 => x"86c72d86",
   977 => x"c72d86c7",
   978 => x"2d86c72d",
   979 => x"86c72d86",
   980 => x"c72d86c7",
   981 => x"2d86c72d",
   982 => x"86c72d86",
   983 => x"c72d86c7",
   984 => x"2d86c72d",
   985 => x"86c72d86",
   986 => x"c72d86c7",
   987 => x"2d86c72d",
   988 => x"86c72d86",
   989 => x"c72d86c7",
   990 => x"2d86c72d",
   991 => x"86c72d86",
   992 => x"c72d86c7",
   993 => x"2d86c72d",
   994 => x"86c72d86",
   995 => x"c72d86c7",
   996 => x"2d86c72d",
   997 => x"86c72d86",
   998 => x"c72d86c7",
   999 => x"2d86c72d",
  1000 => x"86c72d86",
  1001 => x"c72d86c7",
  1002 => x"2d86c72d",
  1003 => x"86c72d86",
  1004 => x"c72d86c7",
  1005 => x"2d86c72d",
  1006 => x"86c72d86",
  1007 => x"c72d86c7",
  1008 => x"2d86c72d",
  1009 => x"86c72d86",
  1010 => x"c72d86c7",
  1011 => x"2d86c72d",
  1012 => x"86c72d86",
  1013 => x"c72d86c7",
  1014 => x"2d86c72d",
  1015 => x"86c72d86",
  1016 => x"c72d86c7",
  1017 => x"2d86c72d",
  1018 => x"86c72d86",
  1019 => x"c72d86c7",
  1020 => x"2d86c72d",
  1021 => x"86c72d86",
  1022 => x"c72d86c7",
  1023 => x"2d86c72d",
  1024 => x"86c72d86",
  1025 => x"c72d86c7",
  1026 => x"2d86c72d",
  1027 => x"86c72d86",
  1028 => x"c72d86c7",
  1029 => x"2d86c72d",
  1030 => x"86c72d86",
  1031 => x"c72d86c7",
  1032 => x"2d86c72d",
  1033 => x"86c72d86",
  1034 => x"c72d86c7",
  1035 => x"2d86c72d",
  1036 => x"86c72d86",
  1037 => x"c72d86c7",
  1038 => x"2d86c72d",
  1039 => x"86c72d86",
  1040 => x"c72d86c7",
  1041 => x"2d86c72d",
  1042 => x"86c72d86",
  1043 => x"c72d86c7",
  1044 => x"2d86c72d",
  1045 => x"86c72d86",
  1046 => x"c72d86c7",
  1047 => x"2d86c72d",
  1048 => x"86c72d86",
  1049 => x"c72d86c7",
  1050 => x"2d86c72d",
  1051 => x"86c72d86",
  1052 => x"c72d86c7",
  1053 => x"2d86c72d",
  1054 => x"86c72d86",
  1055 => x"c72d86c7",
  1056 => x"2d86c72d",
  1057 => x"86c72d86",
  1058 => x"c72d86c7",
  1059 => x"2d86c72d",
  1060 => x"86c72d86",
  1061 => x"c72d86c7",
  1062 => x"2d86c72d",
  1063 => x"86c72d86",
  1064 => x"c72d86c7",
  1065 => x"2d86c72d",
  1066 => x"86c72d86",
  1067 => x"c72d86c7",
  1068 => x"2d86c72d",
  1069 => x"86c72d86",
  1070 => x"c72d86c7",
  1071 => x"2d86c72d",
  1072 => x"86c72d86",
  1073 => x"c72d86c7",
  1074 => x"2d86c72d",
  1075 => x"86c72d86",
  1076 => x"c72d86c7",
  1077 => x"2d86c72d",
  1078 => x"86c72d86",
  1079 => x"c72d86c7",
  1080 => x"2d86c72d",
  1081 => x"86c72d86",
  1082 => x"c72d86c7",
  1083 => x"2d86c72d",
  1084 => x"86c72d86",
  1085 => x"c72d86c7",
  1086 => x"2d86c72d",
  1087 => x"86c72d86",
  1088 => x"c72d86c7",
  1089 => x"2d86c72d",
  1090 => x"82710c02",
  1091 => x"84050d04",
  1092 => x"a00bec0c",
  1093 => x"86c72d86",
  1094 => x"c72d86c7",
  1095 => x"2d86c72d",
  1096 => x"86c72d86",
  1097 => x"c72d86c7",
  1098 => x"2d86c72d",
  1099 => x"86c72d86",
  1100 => x"c72d86c7",
  1101 => x"2d86c72d",
  1102 => x"86c72d86",
  1103 => x"c72d86c7",
  1104 => x"2d86c72d",
  1105 => x"86c72d86",
  1106 => x"c72d86c7",
  1107 => x"2d86c72d",
  1108 => x"86c72d86",
  1109 => x"c72d86c7",
  1110 => x"2d86c72d",
  1111 => x"86c72d86",
  1112 => x"c72d86c7",
  1113 => x"2d86c72d",
  1114 => x"86c72d86",
  1115 => x"c72d86c7",
  1116 => x"2d86c72d",
  1117 => x"86c72d86",
  1118 => x"c72d86c7",
  1119 => x"2d86c72d",
  1120 => x"86c72d86",
  1121 => x"c72d86c7",
  1122 => x"2d86c72d",
  1123 => x"86c72d86",
  1124 => x"c72d86c7",
  1125 => x"2d86c72d",
  1126 => x"86c72d86",
  1127 => x"c72d86c7",
  1128 => x"2d86c72d",
  1129 => x"86c72d86",
  1130 => x"c72d86c7",
  1131 => x"2d86c72d",
  1132 => x"86c72d86",
  1133 => x"c72d86c7",
  1134 => x"2d86c72d",
  1135 => x"86c72d86",
  1136 => x"c72d86c7",
  1137 => x"2d86c72d",
  1138 => x"86c72d86",
  1139 => x"c72d86c7",
  1140 => x"2d86c72d",
  1141 => x"86c72d86",
  1142 => x"c72d86c7",
  1143 => x"2d86c72d",
  1144 => x"86c72d86",
  1145 => x"c72d86c7",
  1146 => x"2d86c72d",
  1147 => x"86c72d86",
  1148 => x"c72d86c7",
  1149 => x"2d86c72d",
  1150 => x"86c72d86",
  1151 => x"c72d86c7",
  1152 => x"2d86c72d",
  1153 => x"86c72d86",
  1154 => x"c72d86c7",
  1155 => x"2d86c72d",
  1156 => x"86c72d86",
  1157 => x"c72d86c7",
  1158 => x"2d86c72d",
  1159 => x"86c72d86",
  1160 => x"c72d86c7",
  1161 => x"2d86c72d",
  1162 => x"86c72d86",
  1163 => x"c72d86c7",
  1164 => x"2d86c72d",
  1165 => x"86c72d86",
  1166 => x"c72d86c7",
  1167 => x"2d86c72d",
  1168 => x"86c72d86",
  1169 => x"c72d86c7",
  1170 => x"2d86c72d",
  1171 => x"86c72d86",
  1172 => x"c72d86c7",
  1173 => x"2d86c72d",
  1174 => x"86c72d86",
  1175 => x"c72d86c7",
  1176 => x"2d86c72d",
  1177 => x"86c72d86",
  1178 => x"c72d86c7",
  1179 => x"2d86c72d",
  1180 => x"86c72d86",
  1181 => x"c72d86c7",
  1182 => x"2d86c72d",
  1183 => x"86c72d86",
  1184 => x"c72d86c7",
  1185 => x"2d86c72d",
  1186 => x"86c72d86",
  1187 => x"c72d86c7",
  1188 => x"2d86c72d",
  1189 => x"86c72d86",
  1190 => x"c72d86c7",
  1191 => x"2d86c72d",
  1192 => x"86c72d86",
  1193 => x"c72d86c7",
  1194 => x"2d86c72d",
  1195 => x"86c72d86",
  1196 => x"c72d86c7",
  1197 => x"2d86c72d",
  1198 => x"86c72d86",
  1199 => x"c72d86c7",
  1200 => x"2d86c72d",
  1201 => x"86c72d86",
  1202 => x"c72d86c7",
  1203 => x"2d86c72d",
  1204 => x"86c72d86",
  1205 => x"c72d86c7",
  1206 => x"2d86c72d",
  1207 => x"86c72d86",
  1208 => x"c72d86c7",
  1209 => x"2d86c72d",
  1210 => x"86c72d86",
  1211 => x"c72d86c7",
  1212 => x"2d86c72d",
  1213 => x"86c72d86",
  1214 => x"c72d86c7",
  1215 => x"2d86c72d",
  1216 => x"86c72d86",
  1217 => x"c72d86c7",
  1218 => x"2d86c72d",
  1219 => x"86c72d86",
  1220 => x"c72d86c7",
  1221 => x"2d86c72d",
  1222 => x"86c72d86",
  1223 => x"c72d86c7",
  1224 => x"2d86c72d",
  1225 => x"86c72d86",
  1226 => x"c72d86c7",
  1227 => x"2d86c72d",
  1228 => x"86c72d86",
  1229 => x"c72d86c7",
  1230 => x"2d86c72d",
  1231 => x"86c72d86",
  1232 => x"c72d86c7",
  1233 => x"2d86c72d",
  1234 => x"86c72d86",
  1235 => x"c72d86c7",
  1236 => x"2d86c72d",
  1237 => x"86c72d86",
  1238 => x"c72d86c7",
  1239 => x"2d86c72d",
  1240 => x"86c72d86",
  1241 => x"c72d86c7",
  1242 => x"2d86c72d",
  1243 => x"86c72d86",
  1244 => x"c72d86c7",
  1245 => x"2d86c72d",
  1246 => x"86c72d86",
  1247 => x"c72d86c7",
  1248 => x"2d86c72d",
  1249 => x"86c72d86",
  1250 => x"c72d86c7",
  1251 => x"2d86c72d",
  1252 => x"86c72d86",
  1253 => x"c72d86c7",
  1254 => x"2d86c72d",
  1255 => x"86c72d86",
  1256 => x"c72d86c7",
  1257 => x"2d86c72d",
  1258 => x"86c72d86",
  1259 => x"c72d86c7",
  1260 => x"2d86c72d",
  1261 => x"86c72d86",
  1262 => x"c72d86c7",
  1263 => x"2d86c72d",
  1264 => x"86c72d86",
  1265 => x"c72d86c7",
  1266 => x"2d86c72d",
  1267 => x"86c72d86",
  1268 => x"c72d86c7",
  1269 => x"2d86c72d",
  1270 => x"86c72d86",
  1271 => x"c72d86c7",
  1272 => x"2d86c72d",
  1273 => x"86c72d86",
  1274 => x"c72d86c7",
  1275 => x"2d86c72d",
  1276 => x"86c72d86",
  1277 => x"c72d86c7",
  1278 => x"2d86c72d",
  1279 => x"86c72d86",
  1280 => x"c72d86c7",
  1281 => x"2d86c72d",
  1282 => x"86c72d86",
  1283 => x"c72d86c7",
  1284 => x"2d86c72d",
  1285 => x"86c72d86",
  1286 => x"c72d86c7",
  1287 => x"2d86c72d",
  1288 => x"86c72d86",
  1289 => x"c72d86c7",
  1290 => x"2d86c72d",
  1291 => x"86c72d86",
  1292 => x"c72d86c7",
  1293 => x"2d86c72d",
  1294 => x"86c72d86",
  1295 => x"c72d86c7",
  1296 => x"2d86c72d",
  1297 => x"86c72d86",
  1298 => x"c72d86c7",
  1299 => x"2d86c72d",
  1300 => x"86c72d86",
  1301 => x"c72d86c7",
  1302 => x"2d86c72d",
  1303 => x"86c72d86",
  1304 => x"c72d86c7",
  1305 => x"2d86c72d",
  1306 => x"86c72d86",
  1307 => x"c72d86c7",
  1308 => x"2d86c72d",
  1309 => x"86c72d86",
  1310 => x"c72d86c7",
  1311 => x"2d86c72d",
  1312 => x"86c72d86",
  1313 => x"c72d86c7",
  1314 => x"2d86c72d",
  1315 => x"86c72d86",
  1316 => x"c72d86c7",
  1317 => x"2d86c72d",
  1318 => x"86c72d86",
  1319 => x"c72d86c7",
  1320 => x"2d86c72d",
  1321 => x"86c72d86",
  1322 => x"c72d86c7",
  1323 => x"2d86c72d",
  1324 => x"86c72d86",
  1325 => x"c72d86c7",
  1326 => x"2d86c72d",
  1327 => x"86c72d86",
  1328 => x"c72d86c7",
  1329 => x"2d86c72d",
  1330 => x"86c72d86",
  1331 => x"c72d86c7",
  1332 => x"2d86c72d",
  1333 => x"86c72d86",
  1334 => x"c72d86c7",
  1335 => x"2d86c72d",
  1336 => x"86c72d86",
  1337 => x"c72d86c7",
  1338 => x"2d86c72d",
  1339 => x"86c72d86",
  1340 => x"c72d86c7",
  1341 => x"2d86c72d",
  1342 => x"86c72d86",
  1343 => x"c72d86c7",
  1344 => x"2d86c72d",
  1345 => x"86c72d86",
  1346 => x"c72d86c7",
  1347 => x"2d86c72d",
  1348 => x"86c72d86",
  1349 => x"c72d86c7",
  1350 => x"2d86c72d",
  1351 => x"86c72d86",
  1352 => x"c72d86c7",
  1353 => x"2d86c72d",
  1354 => x"86c72d86",
  1355 => x"c72d86c7",
  1356 => x"2d86c72d",
  1357 => x"86c72d86",
  1358 => x"c72d86c7",
  1359 => x"2d86c72d",
  1360 => x"86c72d86",
  1361 => x"c72d86c7",
  1362 => x"2d86c72d",
  1363 => x"86c72d86",
  1364 => x"c72d86c7",
  1365 => x"2d86c72d",
  1366 => x"86c72d86",
  1367 => x"c72d86c7",
  1368 => x"2d86c72d",
  1369 => x"86c72d86",
  1370 => x"c72d86c7",
  1371 => x"2d86c72d",
  1372 => x"86c72d86",
  1373 => x"c72d86c7",
  1374 => x"2d86c72d",
  1375 => x"86c72d86",
  1376 => x"c72d86c7",
  1377 => x"2d86c72d",
  1378 => x"86c72d86",
  1379 => x"c72d86c7",
  1380 => x"2d86c72d",
  1381 => x"86c72d86",
  1382 => x"c72d86c7",
  1383 => x"2d86c72d",
  1384 => x"86c72d86",
  1385 => x"c72d86c7",
  1386 => x"2d86c72d",
  1387 => x"86c72d86",
  1388 => x"c72d86c7",
  1389 => x"2d86c72d",
  1390 => x"86c72d86",
  1391 => x"c72d86c7",
  1392 => x"2d86c72d",
  1393 => x"86c72d86",
  1394 => x"c72d86c7",
  1395 => x"2d86c72d",
  1396 => x"86c72d86",
  1397 => x"c72d86c7",
  1398 => x"2d86c72d",
  1399 => x"86c72d86",
  1400 => x"c72d86c7",
  1401 => x"2d86c72d",
  1402 => x"86c72d86",
  1403 => x"c72d86c7",
  1404 => x"2d86c72d",
  1405 => x"86c72d86",
  1406 => x"c72d86c7",
  1407 => x"2d86c72d",
  1408 => x"86c72d86",
  1409 => x"c72d86c7",
  1410 => x"2d86c72d",
  1411 => x"86c72d86",
  1412 => x"c72d86c7",
  1413 => x"2d86c72d",
  1414 => x"86c72d86",
  1415 => x"c72d86c7",
  1416 => x"2d86c72d",
  1417 => x"86c72d86",
  1418 => x"c72d86c7",
  1419 => x"2d86c72d",
  1420 => x"86c72d86",
  1421 => x"c72d86c7",
  1422 => x"2d86c72d",
  1423 => x"86c72d86",
  1424 => x"c72d86c7",
  1425 => x"2d86c72d",
  1426 => x"86c72d86",
  1427 => x"c72d86c7",
  1428 => x"2d86c72d",
  1429 => x"86c72d86",
  1430 => x"c72d86c7",
  1431 => x"2d86c72d",
  1432 => x"86c72d86",
  1433 => x"c72d86c7",
  1434 => x"2d86c72d",
  1435 => x"86c72d86",
  1436 => x"c72d86c7",
  1437 => x"2d86c72d",
  1438 => x"86c72d86",
  1439 => x"c72d86c7",
  1440 => x"2d86c72d",
  1441 => x"86c72d86",
  1442 => x"c72d86c7",
  1443 => x"2d86c72d",
  1444 => x"86c72d86",
  1445 => x"c72d86c7",
  1446 => x"2d86c72d",
  1447 => x"86c72d86",
  1448 => x"c72d86c7",
  1449 => x"2d86c72d",
  1450 => x"86c72d86",
  1451 => x"c72d86c7",
  1452 => x"2d86c72d",
  1453 => x"86c72d86",
  1454 => x"c72d86c7",
  1455 => x"2d86c72d",
  1456 => x"86c72d86",
  1457 => x"c72d86c7",
  1458 => x"2d86c72d",
  1459 => x"86c72d86",
  1460 => x"c72d86c7",
  1461 => x"2d86c72d",
  1462 => x"86c72d86",
  1463 => x"c72d86c7",
  1464 => x"2d86c72d",
  1465 => x"86c72d86",
  1466 => x"c72d86c7",
  1467 => x"2d86c72d",
  1468 => x"86c72d86",
  1469 => x"c72d86c7",
  1470 => x"2d86c72d",
  1471 => x"86c72d86",
  1472 => x"c72d86c7",
  1473 => x"2d86c72d",
  1474 => x"86c72d86",
  1475 => x"c72d86c7",
  1476 => x"2d86c72d",
  1477 => x"86c72d86",
  1478 => x"c72d86c7",
  1479 => x"2d86c72d",
  1480 => x"86c72d86",
  1481 => x"c72d86c7",
  1482 => x"2d86c72d",
  1483 => x"86c72d86",
  1484 => x"c72d86c7",
  1485 => x"2d86c72d",
  1486 => x"86c72d86",
  1487 => x"c72d86c7",
  1488 => x"2d86c72d",
  1489 => x"86c72d86",
  1490 => x"c72d86c7",
  1491 => x"2d86c72d",
  1492 => x"86c72d86",
  1493 => x"c72d86c7",
  1494 => x"2d86c72d",
  1495 => x"86c72d86",
  1496 => x"c72d86c7",
  1497 => x"2d86c72d",
  1498 => x"86c72d86",
  1499 => x"c72d86c7",
  1500 => x"2d86c72d",
  1501 => x"86c72d86",
  1502 => x"c72d86c7",
  1503 => x"2d86c72d",
  1504 => x"86c72d86",
  1505 => x"c72d86c7",
  1506 => x"2d86c72d",
  1507 => x"86c72d86",
  1508 => x"c72d86c7",
  1509 => x"2d86c72d",
  1510 => x"86c72d86",
  1511 => x"c72d86c7",
  1512 => x"2d86c72d",
  1513 => x"86c72d86",
  1514 => x"c72d86c7",
  1515 => x"2d86c72d",
  1516 => x"86c72d86",
  1517 => x"c72d86c7",
  1518 => x"2d86c72d",
  1519 => x"86c72d86",
  1520 => x"c72d86c7",
  1521 => x"2d86c72d",
  1522 => x"86c72d86",
  1523 => x"c72d86c7",
  1524 => x"2d86c72d",
  1525 => x"0402dc05",
  1526 => x"0d8059a2",
  1527 => x"902d810b",
  1528 => x"ec0c7a52",
  1529 => x"80e6a851",
  1530 => x"80d6952d",
  1531 => x"80e68c08",
  1532 => x"792e80f7",
  1533 => x"3880e6ac",
  1534 => x"0870f80c",
  1535 => x"79ff1256",
  1536 => x"59557379",
  1537 => x"2e8b3881",
  1538 => x"1874812a",
  1539 => x"555873f7",
  1540 => x"38f71858",
  1541 => x"81598075",
  1542 => x"2580d038",
  1543 => x"77527351",
  1544 => x"84a82d80",
  1545 => x"e7805280",
  1546 => x"e6a85180",
  1547 => x"d8eb2d80",
  1548 => x"e68c0880",
  1549 => x"2e9b3880",
  1550 => x"e7805783",
  1551 => x"fc567670",
  1552 => x"84055808",
  1553 => x"e80cfc16",
  1554 => x"56758025",
  1555 => x"f138b0d9",
  1556 => x"0480e68c",
  1557 => x"08598480",
  1558 => x"5580e6a8",
  1559 => x"5180d8ba",
  1560 => x"2dfc8015",
  1561 => x"81155555",
  1562 => x"b0960484",
  1563 => x"0bec0c78",
  1564 => x"802e8e38",
  1565 => x"80e2e451",
  1566 => x"b98b2db7",
  1567 => x"8b2db188",
  1568 => x"0480e3dc",
  1569 => x"51b98b2d",
  1570 => x"7880e68c",
  1571 => x"0c02a405",
  1572 => x"0d0402f4",
  1573 => x"050d840b",
  1574 => x"ec0cb6be",
  1575 => x"2db2ec2d",
  1576 => x"81f92d83",
  1577 => x"52b6a12d",
  1578 => x"8151858d",
  1579 => x"2dff1252",
  1580 => x"718025f1",
  1581 => x"38840bec",
  1582 => x"0c80e0f4",
  1583 => x"5186a02d",
  1584 => x"80ccb52d",
  1585 => x"80e68c08",
  1586 => x"802e8189",
  1587 => x"3880e18c",
  1588 => x"5186a02d",
  1589 => x"800bf00c",
  1590 => x"80e1a051",
  1591 => x"afd52d81",
  1592 => x"0bf00caf",
  1593 => x"d55180df",
  1594 => x"c22d80e2",
  1595 => x"e451b98b",
  1596 => x"2db6f72d",
  1597 => x"b2f82db9",
  1598 => x"9e2d800b",
  1599 => x"80e2f80b",
  1600 => x"80f52d53",
  1601 => x"5371732e",
  1602 => x"83388453",
  1603 => x"80e3840b",
  1604 => x"80f52d52",
  1605 => x"71802e85",
  1606 => x"38728807",
  1607 => x"5380e390",
  1608 => x"0b80f52d",
  1609 => x"5271802e",
  1610 => x"85387290",
  1611 => x"075380e4",
  1612 => x"c808852a",
  1613 => x"70810651",
  1614 => x"5271802e",
  1615 => x"853872a0",
  1616 => x"075372fc",
  1617 => x"0c865280",
  1618 => x"e68c0883",
  1619 => x"38845271",
  1620 => x"ec0cb1f4",
  1621 => x"04800b80",
  1622 => x"e68c0c02",
  1623 => x"8c050d04",
  1624 => x"71980c04",
  1625 => x"ffb00880",
  1626 => x"e68c0c04",
  1627 => x"810bffb0",
  1628 => x"0c04800b",
  1629 => x"ffb00c04",
  1630 => x"02f4050d",
  1631 => x"80e6b451",
  1632 => x"b58b2dff",
  1633 => x"0b80e68c",
  1634 => x"08258188",
  1635 => x"3880e68c",
  1636 => x"0881f02e",
  1637 => x"0981068a",
  1638 => x"38810b80",
  1639 => x"e4c00cb4",
  1640 => x"940480e6",
  1641 => x"8c0881e0",
  1642 => x"2e098106",
  1643 => x"8a38810b",
  1644 => x"80e4c40c",
  1645 => x"b4940480",
  1646 => x"e68c0852",
  1647 => x"80e4c408",
  1648 => x"802e8938",
  1649 => x"80e68c08",
  1650 => x"81800552",
  1651 => x"71842c72",
  1652 => x"8f065353",
  1653 => x"80e4c008",
  1654 => x"802e9a38",
  1655 => x"72842980",
  1656 => x"e4800572",
  1657 => x"1381712b",
  1658 => x"70097308",
  1659 => x"06730c51",
  1660 => x"5353b488",
  1661 => x"04728429",
  1662 => x"80e48005",
  1663 => x"72138371",
  1664 => x"2b720807",
  1665 => x"720c5353",
  1666 => x"800b80e4",
  1667 => x"c40c800b",
  1668 => x"80e4c00c",
  1669 => x"800b80e6",
  1670 => x"8c0c028c",
  1671 => x"050d0402",
  1672 => x"f8050d80",
  1673 => x"e480528f",
  1674 => x"51807270",
  1675 => x"8405540c",
  1676 => x"ff115170",
  1677 => x"8025f238",
  1678 => x"0288050d",
  1679 => x"0402f005",
  1680 => x"0d7551b2",
  1681 => x"f22d7082",
  1682 => x"2cfc0680",
  1683 => x"e4801172",
  1684 => x"109e0671",
  1685 => x"0870722a",
  1686 => x"70830682",
  1687 => x"742b7009",
  1688 => x"7406760c",
  1689 => x"54515657",
  1690 => x"535153b2",
  1691 => x"ec2d7180",
  1692 => x"e68c0c02",
  1693 => x"90050d04",
  1694 => x"02fc050d",
  1695 => x"72518071",
  1696 => x"0c800b84",
  1697 => x"120c0284",
  1698 => x"050d0402",
  1699 => x"f0050d75",
  1700 => x"70088412",
  1701 => x"08535353",
  1702 => x"ff547171",
  1703 => x"2ea838b2",
  1704 => x"f22d8413",
  1705 => x"08708429",
  1706 => x"14881170",
  1707 => x"087081ff",
  1708 => x"06841808",
  1709 => x"81118706",
  1710 => x"841a0c53",
  1711 => x"51555151",
  1712 => x"51b2ec2d",
  1713 => x"71547380",
  1714 => x"e68c0c02",
  1715 => x"90050d04",
  1716 => x"02f4050d",
  1717 => x"b2f22de0",
  1718 => x"08708b2a",
  1719 => x"70810651",
  1720 => x"52537080",
  1721 => x"2ea13880",
  1722 => x"e6b40870",
  1723 => x"842980e6",
  1724 => x"bc057481",
  1725 => x"ff06710c",
  1726 => x"515180e6",
  1727 => x"b4088111",
  1728 => x"870680e6",
  1729 => x"b40c5172",
  1730 => x"8c2cbf06",
  1731 => x"80e6dc0c",
  1732 => x"800b80e6",
  1733 => x"e00cb2e4",
  1734 => x"2db2ec2d",
  1735 => x"028c050d",
  1736 => x"0402fc05",
  1737 => x"0db2f22d",
  1738 => x"810b80e6",
  1739 => x"e00cb2ec",
  1740 => x"2d80e6e0",
  1741 => x"085170f9",
  1742 => x"38028405",
  1743 => x"0d0402fc",
  1744 => x"050d80e6",
  1745 => x"b451b4f8",
  1746 => x"2db49f2d",
  1747 => x"b5d051b2",
  1748 => x"e02d0284",
  1749 => x"050d0402",
  1750 => x"fc050d8f",
  1751 => x"cf5186c7",
  1752 => x"2dff1151",
  1753 => x"708025f6",
  1754 => x"38028405",
  1755 => x"0d0480e6",
  1756 => x"ec0880e6",
  1757 => x"8c0c0402",
  1758 => x"fc050d81",
  1759 => x"0b80e4cc",
  1760 => x"0c815185",
  1761 => x"8d2d0284",
  1762 => x"050d0402",
  1763 => x"fc050db7",
  1764 => x"9504b2f8",
  1765 => x"2d8751b4",
  1766 => x"bd2d80e6",
  1767 => x"8c08f338",
  1768 => x"80e68c08",
  1769 => x"80e4cc0c",
  1770 => x"80e68c08",
  1771 => x"51858d2d",
  1772 => x"0284050d",
  1773 => x"0402ec05",
  1774 => x"0d765480",
  1775 => x"52870b88",
  1776 => x"1580f52d",
  1777 => x"56537472",
  1778 => x"248338a0",
  1779 => x"53725183",
  1780 => x"842d8112",
  1781 => x"8b1580f5",
  1782 => x"2d545272",
  1783 => x"7225de38",
  1784 => x"0294050d",
  1785 => x"0402f005",
  1786 => x"0d80e6ec",
  1787 => x"085481f9",
  1788 => x"2d800b80",
  1789 => x"e6f00c73",
  1790 => x"08802e81",
  1791 => x"8938820b",
  1792 => x"80e6a00c",
  1793 => x"80e6f008",
  1794 => x"8f0680e6",
  1795 => x"9c0c7308",
  1796 => x"5271832e",
  1797 => x"96387183",
  1798 => x"26893871",
  1799 => x"812eb038",
  1800 => x"b8ef0471",
  1801 => x"852ea038",
  1802 => x"b8ef0488",
  1803 => x"1480f52d",
  1804 => x"84150880",
  1805 => x"e1ac5354",
  1806 => x"5286a02d",
  1807 => x"71842913",
  1808 => x"70085252",
  1809 => x"b8f30473",
  1810 => x"51b7b52d",
  1811 => x"b8ef0480",
  1812 => x"e4c80888",
  1813 => x"15082c70",
  1814 => x"81065152",
  1815 => x"71802e88",
  1816 => x"3880e1b0",
  1817 => x"51b8ec04",
  1818 => x"80e1b451",
  1819 => x"86a02d84",
  1820 => x"14085186",
  1821 => x"a02d80e6",
  1822 => x"f0088105",
  1823 => x"80e6f00c",
  1824 => x"8c1454b7",
  1825 => x"f7040290",
  1826 => x"050d0471",
  1827 => x"80e6ec0c",
  1828 => x"b7e52d80",
  1829 => x"e6f008ff",
  1830 => x"0580e6f4",
  1831 => x"0c0402e8",
  1832 => x"050d80e6",
  1833 => x"ec0880e6",
  1834 => x"f8085755",
  1835 => x"8751b4bd",
  1836 => x"2d80e68c",
  1837 => x"08812a70",
  1838 => x"81065152",
  1839 => x"71802ea1",
  1840 => x"38b9c704",
  1841 => x"b2f82d87",
  1842 => x"51b4bd2d",
  1843 => x"80e68c08",
  1844 => x"f33880e4",
  1845 => x"cc088132",
  1846 => x"7080e4cc",
  1847 => x"0c51858d",
  1848 => x"2d80e6dc",
  1849 => x"08a00652",
  1850 => x"80722598",
  1851 => x"38b6d72d",
  1852 => x"b2f82d80",
  1853 => x"e4cc0881",
  1854 => x"327080e4",
  1855 => x"cc0c7052",
  1856 => x"52858d2d",
  1857 => x"800b80e6",
  1858 => x"e40c800b",
  1859 => x"80e6e80c",
  1860 => x"80e4cc08",
  1861 => x"83ae3880",
  1862 => x"da51b4bd",
  1863 => x"2d80e68c",
  1864 => x"08802e8c",
  1865 => x"3880e6e4",
  1866 => x"08818007",
  1867 => x"80e6e40c",
  1868 => x"80d951b4",
  1869 => x"bd2d80e6",
  1870 => x"8c08802e",
  1871 => x"8c3880e6",
  1872 => x"e40880c0",
  1873 => x"0780e6e4",
  1874 => x"0c819451",
  1875 => x"b4bd2d80",
  1876 => x"e68c0880",
  1877 => x"2e8b3880",
  1878 => x"e6e40890",
  1879 => x"0780e6e4",
  1880 => x"0c819151",
  1881 => x"b4bd2d80",
  1882 => x"e68c0880",
  1883 => x"2e8b3880",
  1884 => x"e6e408a0",
  1885 => x"0780e6e4",
  1886 => x"0c81f551",
  1887 => x"b4bd2d80",
  1888 => x"e68c0880",
  1889 => x"2e8b3880",
  1890 => x"e6e40881",
  1891 => x"0780e6e4",
  1892 => x"0c81f251",
  1893 => x"b4bd2d80",
  1894 => x"e68c0880",
  1895 => x"2e8b3880",
  1896 => x"e6e40882",
  1897 => x"0780e6e4",
  1898 => x"0c81eb51",
  1899 => x"b4bd2d80",
  1900 => x"e68c0880",
  1901 => x"2e8b3880",
  1902 => x"e6e40884",
  1903 => x"0780e6e4",
  1904 => x"0c81f451",
  1905 => x"b4bd2d80",
  1906 => x"e68c0880",
  1907 => x"2e8b3880",
  1908 => x"e6e40888",
  1909 => x"0780e6e4",
  1910 => x"0c80d851",
  1911 => x"b4bd2d80",
  1912 => x"e68c0880",
  1913 => x"2e8c3880",
  1914 => x"e6e80881",
  1915 => x"800780e6",
  1916 => x"e80c9251",
  1917 => x"b4bd2d80",
  1918 => x"e68c0880",
  1919 => x"2e8c3880",
  1920 => x"e6e80880",
  1921 => x"c00780e6",
  1922 => x"e80c9451",
  1923 => x"b4bd2d80",
  1924 => x"e68c0880",
  1925 => x"2e8b3880",
  1926 => x"e6e80890",
  1927 => x"0780e6e8",
  1928 => x"0c9151b4",
  1929 => x"bd2d80e6",
  1930 => x"8c08802e",
  1931 => x"8b3880e6",
  1932 => x"e808a007",
  1933 => x"80e6e80c",
  1934 => x"9d51b4bd",
  1935 => x"2d80e68c",
  1936 => x"08802e8b",
  1937 => x"3880e6e8",
  1938 => x"08810780",
  1939 => x"e6e80c9b",
  1940 => x"51b4bd2d",
  1941 => x"80e68c08",
  1942 => x"802e8b38",
  1943 => x"80e6e808",
  1944 => x"820780e6",
  1945 => x"e80c9c51",
  1946 => x"b4bd2d80",
  1947 => x"e68c0880",
  1948 => x"2e8b3880",
  1949 => x"e6e80884",
  1950 => x"0780e6e8",
  1951 => x"0ca351b4",
  1952 => x"bd2d80e6",
  1953 => x"8c08802e",
  1954 => x"8b3880e6",
  1955 => x"e8088807",
  1956 => x"80e6e80c",
  1957 => x"9651b4bd",
  1958 => x"2d80e68c",
  1959 => x"08802e84",
  1960 => x"3894bf2d",
  1961 => x"9e51b4bd",
  1962 => x"2d80e68c",
  1963 => x"08802e84",
  1964 => x"3886ee2d",
  1965 => x"81fd51b4",
  1966 => x"bd2d81fa",
  1967 => x"51b4bd2d",
  1968 => x"80c3ee04",
  1969 => x"81f551b4",
  1970 => x"bd2d80e6",
  1971 => x"8c08812a",
  1972 => x"70810651",
  1973 => x"52718e38",
  1974 => x"80e6dc08",
  1975 => x"90065280",
  1976 => x"722580c2",
  1977 => x"3880e6dc",
  1978 => x"08900652",
  1979 => x"80722584",
  1980 => x"38b6d72d",
  1981 => x"80e6f408",
  1982 => x"5271802e",
  1983 => x"8a38ff12",
  1984 => x"80e6f40c",
  1985 => x"bea60480",
  1986 => x"e6f00810",
  1987 => x"80e6f008",
  1988 => x"05708429",
  1989 => x"16515288",
  1990 => x"1208802e",
  1991 => x"8938ff51",
  1992 => x"88120852",
  1993 => x"712d81f2",
  1994 => x"51b4bd2d",
  1995 => x"80e68c08",
  1996 => x"812a7081",
  1997 => x"06515271",
  1998 => x"8e3880e6",
  1999 => x"dc088806",
  2000 => x"52807225",
  2001 => x"80c33880",
  2002 => x"e6dc0888",
  2003 => x"06528072",
  2004 => x"258438b6",
  2005 => x"d72d80e6",
  2006 => x"f008ff11",
  2007 => x"80e6f408",
  2008 => x"56535373",
  2009 => x"72258a38",
  2010 => x"811480e6",
  2011 => x"f40cbf89",
  2012 => x"04721013",
  2013 => x"70842916",
  2014 => x"51528812",
  2015 => x"08802e89",
  2016 => x"38fe5188",
  2017 => x"12085271",
  2018 => x"2d81fd51",
  2019 => x"b4bd2d80",
  2020 => x"e68c0881",
  2021 => x"2a708106",
  2022 => x"51527180",
  2023 => x"2eb13880",
  2024 => x"e6f40880",
  2025 => x"2e8a3880",
  2026 => x"0b80e6f4",
  2027 => x"0cbfcf04",
  2028 => x"80e6f008",
  2029 => x"1080e6f0",
  2030 => x"08057084",
  2031 => x"29165152",
  2032 => x"88120880",
  2033 => x"2e8938fd",
  2034 => x"51881208",
  2035 => x"52712d81",
  2036 => x"fa51b4bd",
  2037 => x"2d80e68c",
  2038 => x"08812a70",
  2039 => x"81065152",
  2040 => x"71802eb2",
  2041 => x"3880e6f0",
  2042 => x"08ff1154",
  2043 => x"5280e6f4",
  2044 => x"0873258a",
  2045 => x"387280e6",
  2046 => x"f40c80c0",
  2047 => x"96047110",
  2048 => x"12708429",
  2049 => x"16515288",
  2050 => x"1208802e",
  2051 => x"8938fc51",
  2052 => x"88120852",
  2053 => x"712d80e6",
  2054 => x"f4087053",
  2055 => x"5473802e",
  2056 => x"8b388c15",
  2057 => x"ff155555",
  2058 => x"80c09d04",
  2059 => x"820b80e6",
  2060 => x"a00c718f",
  2061 => x"0680e69c",
  2062 => x"0c81eb51",
  2063 => x"b4bd2d80",
  2064 => x"e68c0881",
  2065 => x"2a708106",
  2066 => x"51527180",
  2067 => x"2ead3874",
  2068 => x"08852e09",
  2069 => x"8106a438",
  2070 => x"881580f5",
  2071 => x"2dff0552",
  2072 => x"71881681",
  2073 => x"b72d7198",
  2074 => x"2b527180",
  2075 => x"25883880",
  2076 => x"0b881681",
  2077 => x"b72d7451",
  2078 => x"b7b52d81",
  2079 => x"f451b4bd",
  2080 => x"2d80e68c",
  2081 => x"08812a70",
  2082 => x"81065152",
  2083 => x"71802eb3",
  2084 => x"38740885",
  2085 => x"2e098106",
  2086 => x"aa388815",
  2087 => x"80f52d81",
  2088 => x"05527188",
  2089 => x"1681b72d",
  2090 => x"7181ff06",
  2091 => x"8b1680f5",
  2092 => x"2d545272",
  2093 => x"72278738",
  2094 => x"72881681",
  2095 => x"b72d7451",
  2096 => x"b7b52d80",
  2097 => x"da51b4bd",
  2098 => x"2d80e68c",
  2099 => x"08812a70",
  2100 => x"81065152",
  2101 => x"718e3880",
  2102 => x"e6dc0881",
  2103 => x"06528072",
  2104 => x"2581c238",
  2105 => x"80e6ec08",
  2106 => x"80e6dc08",
  2107 => x"81065353",
  2108 => x"80722584",
  2109 => x"38b6d72d",
  2110 => x"80e6f408",
  2111 => x"5473802e",
  2112 => x"8b388c13",
  2113 => x"ff155553",
  2114 => x"80c1fd04",
  2115 => x"72085271",
  2116 => x"822ea838",
  2117 => x"7182268a",
  2118 => x"3871812e",
  2119 => x"ad3880c3",
  2120 => x"a5047183",
  2121 => x"2eb73871",
  2122 => x"842e0981",
  2123 => x"0680f638",
  2124 => x"88130851",
  2125 => x"b98b2d80",
  2126 => x"c3a50480",
  2127 => x"e6f40851",
  2128 => x"88130852",
  2129 => x"712d80c3",
  2130 => x"a504810b",
  2131 => x"8814082b",
  2132 => x"80e4c808",
  2133 => x"3280e4c8",
  2134 => x"0c80c2f8",
  2135 => x"04881380",
  2136 => x"f52d8105",
  2137 => x"8b1480f5",
  2138 => x"2d535471",
  2139 => x"74248338",
  2140 => x"80547388",
  2141 => x"1481b72d",
  2142 => x"b7e52d80",
  2143 => x"c3a50475",
  2144 => x"08802ea4",
  2145 => x"38750851",
  2146 => x"b4bd2d80",
  2147 => x"e68c0881",
  2148 => x"06527180",
  2149 => x"2e8c3880",
  2150 => x"e6f40851",
  2151 => x"84160852",
  2152 => x"712d8816",
  2153 => x"5675d838",
  2154 => x"8054800b",
  2155 => x"80e6a00c",
  2156 => x"738f0680",
  2157 => x"e69c0ca0",
  2158 => x"527380e6",
  2159 => x"f4082e09",
  2160 => x"81069938",
  2161 => x"80e6f008",
  2162 => x"ff057432",
  2163 => x"70098105",
  2164 => x"7072079f",
  2165 => x"2a917131",
  2166 => x"51515353",
  2167 => x"71518384",
  2168 => x"2d811454",
  2169 => x"8e7425c2",
  2170 => x"3880e4cc",
  2171 => x"08527180",
  2172 => x"e68c0c02",
  2173 => x"98050d04",
  2174 => x"02f4050d",
  2175 => x"d45281ff",
  2176 => x"720c7108",
  2177 => x"5381ff72",
  2178 => x"0c72882b",
  2179 => x"83fe8006",
  2180 => x"72087081",
  2181 => x"ff065152",
  2182 => x"5381ff72",
  2183 => x"0c727107",
  2184 => x"882b7208",
  2185 => x"7081ff06",
  2186 => x"51525381",
  2187 => x"ff720c72",
  2188 => x"7107882b",
  2189 => x"72087081",
  2190 => x"ff067207",
  2191 => x"80e68c0c",
  2192 => x"5253028c",
  2193 => x"050d0402",
  2194 => x"f4050d74",
  2195 => x"767181ff",
  2196 => x"06d40c53",
  2197 => x"5380e6fc",
  2198 => x"08853871",
  2199 => x"892b5271",
  2200 => x"982ad40c",
  2201 => x"71902a70",
  2202 => x"81ff06d4",
  2203 => x"0c517188",
  2204 => x"2a7081ff",
  2205 => x"06d40c51",
  2206 => x"7181ff06",
  2207 => x"d40c7290",
  2208 => x"2a7081ff",
  2209 => x"06d40c51",
  2210 => x"d4087081",
  2211 => x"ff065151",
  2212 => x"82b8bf52",
  2213 => x"7081ff2e",
  2214 => x"09810694",
  2215 => x"3881ff0b",
  2216 => x"d40cd408",
  2217 => x"7081ff06",
  2218 => x"ff145451",
  2219 => x"5171e538",
  2220 => x"7080e68c",
  2221 => x"0c028c05",
  2222 => x"0d0402fc",
  2223 => x"050d81c7",
  2224 => x"5181ff0b",
  2225 => x"d40cff11",
  2226 => x"51708025",
  2227 => x"f4380284",
  2228 => x"050d0402",
  2229 => x"f4050d81",
  2230 => x"ff0bd40c",
  2231 => x"93538052",
  2232 => x"87fc80c1",
  2233 => x"5180c4c7",
  2234 => x"2d80e68c",
  2235 => x"088c3881",
  2236 => x"ff0bd40c",
  2237 => x"815380c6",
  2238 => x"840480c5",
  2239 => x"ba2dff13",
  2240 => x"5372db38",
  2241 => x"7280e68c",
  2242 => x"0c028c05",
  2243 => x"0d0402ec",
  2244 => x"050d810b",
  2245 => x"80e6fc0c",
  2246 => x"8454d008",
  2247 => x"708f2a70",
  2248 => x"81065151",
  2249 => x"5372f338",
  2250 => x"72d00c80",
  2251 => x"c5ba2d80",
  2252 => x"e1b85186",
  2253 => x"a02dd008",
  2254 => x"708f2a70",
  2255 => x"81065151",
  2256 => x"5372f338",
  2257 => x"810bd00c",
  2258 => x"b1538052",
  2259 => x"84d480c0",
  2260 => x"5180c4c7",
  2261 => x"2d80e68c",
  2262 => x"08812e94",
  2263 => x"3872822e",
  2264 => x"80c438ff",
  2265 => x"135372e2",
  2266 => x"38ff1454",
  2267 => x"73ffab38",
  2268 => x"80c5ba2d",
  2269 => x"83aa5284",
  2270 => x"9c80c851",
  2271 => x"80c4c72d",
  2272 => x"80e68c08",
  2273 => x"812e0981",
  2274 => x"06943880",
  2275 => x"c3f82d80",
  2276 => x"e68c0883",
  2277 => x"ffff0653",
  2278 => x"7283aa2e",
  2279 => x"a33880c5",
  2280 => x"d32d80c7",
  2281 => x"ba0480e1",
  2282 => x"c45186a0",
  2283 => x"2d805380",
  2284 => x"c9980480",
  2285 => x"e1dc5186",
  2286 => x"a02d8054",
  2287 => x"80c8e804",
  2288 => x"81ff0bd4",
  2289 => x"0cb15480",
  2290 => x"c5ba2d8f",
  2291 => x"cf538052",
  2292 => x"87fc80f7",
  2293 => x"5180c4c7",
  2294 => x"2d80e68c",
  2295 => x"085580e6",
  2296 => x"8c08812e",
  2297 => x"0981069e",
  2298 => x"3881ff0b",
  2299 => x"d40c820a",
  2300 => x"52849c80",
  2301 => x"e95180c4",
  2302 => x"c72d80e6",
  2303 => x"8c08802e",
  2304 => x"8f3880c5",
  2305 => x"ba2dff13",
  2306 => x"5372c338",
  2307 => x"80c8db04",
  2308 => x"81ff0bd4",
  2309 => x"0c80e68c",
  2310 => x"085287fc",
  2311 => x"80fa5180",
  2312 => x"c4c72d80",
  2313 => x"e68c08b3",
  2314 => x"3881ff0b",
  2315 => x"d40cd408",
  2316 => x"5381ff0b",
  2317 => x"d40c81ff",
  2318 => x"0bd40c81",
  2319 => x"ff0bd40c",
  2320 => x"81ff0bd4",
  2321 => x"0c72862a",
  2322 => x"70810676",
  2323 => x"56515372",
  2324 => x"973880e6",
  2325 => x"8c085480",
  2326 => x"c8e80473",
  2327 => x"822efed3",
  2328 => x"38ff1454",
  2329 => x"73fee038",
  2330 => x"7380e6fc",
  2331 => x"0c738c38",
  2332 => x"815287fc",
  2333 => x"80d05180",
  2334 => x"c4c72d81",
  2335 => x"ff0bd40c",
  2336 => x"d008708f",
  2337 => x"2a708106",
  2338 => x"51515372",
  2339 => x"f33872d0",
  2340 => x"0c81ff0b",
  2341 => x"d40c8153",
  2342 => x"7280e68c",
  2343 => x"0c029405",
  2344 => x"0d0402e8",
  2345 => x"050d7855",
  2346 => x"805681ff",
  2347 => x"0bd40cd0",
  2348 => x"08708f2a",
  2349 => x"70810651",
  2350 => x"515372f3",
  2351 => x"3882810b",
  2352 => x"d00c81ff",
  2353 => x"0bd40c77",
  2354 => x"5287fc80",
  2355 => x"d15180c4",
  2356 => x"c72d80db",
  2357 => x"c6df5480",
  2358 => x"e68c0880",
  2359 => x"2e8c3880",
  2360 => x"e1fc5186",
  2361 => x"a02d80ca",
  2362 => x"c00481ff",
  2363 => x"0bd40cd4",
  2364 => x"087081ff",
  2365 => x"06515372",
  2366 => x"81fe2e09",
  2367 => x"8106a038",
  2368 => x"80ff5380",
  2369 => x"c3f82d80",
  2370 => x"e68c0875",
  2371 => x"70840557",
  2372 => x"0cff1353",
  2373 => x"728025eb",
  2374 => x"38815680",
  2375 => x"caa504ff",
  2376 => x"145473c6",
  2377 => x"3881ff0b",
  2378 => x"d40c81ff",
  2379 => x"0bd40cd0",
  2380 => x"08708f2a",
  2381 => x"70810651",
  2382 => x"515372f3",
  2383 => x"3872d00c",
  2384 => x"7580e68c",
  2385 => x"0c029805",
  2386 => x"0d0402e8",
  2387 => x"050d7779",
  2388 => x"7b585555",
  2389 => x"80537276",
  2390 => x"25a53874",
  2391 => x"70810556",
  2392 => x"80f52d74",
  2393 => x"70810556",
  2394 => x"80f52d52",
  2395 => x"5271712e",
  2396 => x"87388151",
  2397 => x"80cb8104",
  2398 => x"81135380",
  2399 => x"cad60480",
  2400 => x"517080e6",
  2401 => x"8c0c0298",
  2402 => x"050d0402",
  2403 => x"ec050d76",
  2404 => x"5574802e",
  2405 => x"80c4389a",
  2406 => x"1580e02d",
  2407 => x"5180d9c6",
  2408 => x"2d80e68c",
  2409 => x"0880e68c",
  2410 => x"0880edb0",
  2411 => x"0c80e68c",
  2412 => x"08545480",
  2413 => x"ed8c0880",
  2414 => x"2e9b3894",
  2415 => x"1580e02d",
  2416 => x"5180d9c6",
  2417 => x"2d80e68c",
  2418 => x"08902b83",
  2419 => x"fff00a06",
  2420 => x"70750751",
  2421 => x"537280ed",
  2422 => x"b00c80ed",
  2423 => x"b0085372",
  2424 => x"802e9e38",
  2425 => x"80ed8408",
  2426 => x"fe147129",
  2427 => x"80ed9808",
  2428 => x"0580edb4",
  2429 => x"0c70842b",
  2430 => x"80ed900c",
  2431 => x"5480ccb0",
  2432 => x"0480ed9c",
  2433 => x"0880edb0",
  2434 => x"0c80eda0",
  2435 => x"0880edb4",
  2436 => x"0c80ed8c",
  2437 => x"08802e8c",
  2438 => x"3880ed84",
  2439 => x"08842b53",
  2440 => x"80ccab04",
  2441 => x"80eda408",
  2442 => x"842b5372",
  2443 => x"80ed900c",
  2444 => x"0294050d",
  2445 => x"0402d805",
  2446 => x"0d800b80",
  2447 => x"ed8c0c84",
  2448 => x"5480c68e",
  2449 => x"2d80e68c",
  2450 => x"08802e99",
  2451 => x"3880e780",
  2452 => x"52805180",
  2453 => x"c9a22d80",
  2454 => x"e68c0880",
  2455 => x"2e8738fe",
  2456 => x"5480cced",
  2457 => x"04ff1454",
  2458 => x"738024d5",
  2459 => x"38738e38",
  2460 => x"80e28c51",
  2461 => x"86a02d73",
  2462 => x"5580d2d1",
  2463 => x"04805681",
  2464 => x"0b80edb8",
  2465 => x"0c885380",
  2466 => x"e2a05280",
  2467 => x"e7b65180",
  2468 => x"caca2d80",
  2469 => x"e68c0876",
  2470 => x"2e098106",
  2471 => x"893880e6",
  2472 => x"8c0880ed",
  2473 => x"b80c8853",
  2474 => x"80e2ac52",
  2475 => x"80e7d251",
  2476 => x"80caca2d",
  2477 => x"80e68c08",
  2478 => x"893880e6",
  2479 => x"8c0880ed",
  2480 => x"b80c80ed",
  2481 => x"b808802e",
  2482 => x"81853880",
  2483 => x"eac60b80",
  2484 => x"f52d80ea",
  2485 => x"c70b80f5",
  2486 => x"2d71982b",
  2487 => x"71902b07",
  2488 => x"80eac80b",
  2489 => x"80f52d70",
  2490 => x"882b7207",
  2491 => x"80eac90b",
  2492 => x"80f52d71",
  2493 => x"0780eafe",
  2494 => x"0b80f52d",
  2495 => x"80eaff0b",
  2496 => x"80f52d71",
  2497 => x"882b0753",
  2498 => x"5f54525a",
  2499 => x"56575573",
  2500 => x"81abaa2e",
  2501 => x"09810690",
  2502 => x"38755180",
  2503 => x"d9952d80",
  2504 => x"e68c0856",
  2505 => x"80ceb704",
  2506 => x"7382d4d5",
  2507 => x"2e893880",
  2508 => x"e2b85180",
  2509 => x"cf870480",
  2510 => x"e7805275",
  2511 => x"5180c9a2",
  2512 => x"2d80e68c",
  2513 => x"085580e6",
  2514 => x"8c08802e",
  2515 => x"84833888",
  2516 => x"5380e2ac",
  2517 => x"5280e7d2",
  2518 => x"5180caca",
  2519 => x"2d80e68c",
  2520 => x"088b3881",
  2521 => x"0b80ed8c",
  2522 => x"0c80cf8e",
  2523 => x"04885380",
  2524 => x"e2a05280",
  2525 => x"e7b65180",
  2526 => x"caca2d80",
  2527 => x"e68c0880",
  2528 => x"2e8c3880",
  2529 => x"e2cc5186",
  2530 => x"a02d80cf",
  2531 => x"ed0480ea",
  2532 => x"fe0b80f5",
  2533 => x"2d547380",
  2534 => x"d52e0981",
  2535 => x"0680ce38",
  2536 => x"80eaff0b",
  2537 => x"80f52d54",
  2538 => x"7381aa2e",
  2539 => x"098106bd",
  2540 => x"38800b80",
  2541 => x"e7800b80",
  2542 => x"f52d5654",
  2543 => x"7481e92e",
  2544 => x"83388154",
  2545 => x"7481eb2e",
  2546 => x"8c388055",
  2547 => x"73752e09",
  2548 => x"810682fd",
  2549 => x"3880e78b",
  2550 => x"0b80f52d",
  2551 => x"55748e38",
  2552 => x"80e78c0b",
  2553 => x"80f52d54",
  2554 => x"73822e87",
  2555 => x"38805580",
  2556 => x"d2d10480",
  2557 => x"e78d0b80",
  2558 => x"f52d7080",
  2559 => x"ed840cff",
  2560 => x"0580ed88",
  2561 => x"0c80e78e",
  2562 => x"0b80f52d",
  2563 => x"80e78f0b",
  2564 => x"80f52d58",
  2565 => x"76057782",
  2566 => x"80290570",
  2567 => x"80ed940c",
  2568 => x"80e7900b",
  2569 => x"80f52d70",
  2570 => x"80eda80c",
  2571 => x"80ed8c08",
  2572 => x"59575876",
  2573 => x"802e81b9",
  2574 => x"38885380",
  2575 => x"e2ac5280",
  2576 => x"e7d25180",
  2577 => x"caca2d80",
  2578 => x"e68c0882",
  2579 => x"843880ed",
  2580 => x"84087084",
  2581 => x"2b80ed90",
  2582 => x"0c7080ed",
  2583 => x"a40c80e7",
  2584 => x"a50b80f5",
  2585 => x"2d80e7a4",
  2586 => x"0b80f52d",
  2587 => x"71828029",
  2588 => x"0580e7a6",
  2589 => x"0b80f52d",
  2590 => x"70848080",
  2591 => x"291280e7",
  2592 => x"a70b80f5",
  2593 => x"2d708180",
  2594 => x"0a291270",
  2595 => x"80edac0c",
  2596 => x"80eda808",
  2597 => x"712980ed",
  2598 => x"94080570",
  2599 => x"80ed980c",
  2600 => x"80e7ad0b",
  2601 => x"80f52d80",
  2602 => x"e7ac0b80",
  2603 => x"f52d7182",
  2604 => x"80290580",
  2605 => x"e7ae0b80",
  2606 => x"f52d7084",
  2607 => x"80802912",
  2608 => x"80e7af0b",
  2609 => x"80f52d70",
  2610 => x"982b81f0",
  2611 => x"0a067205",
  2612 => x"7080ed9c",
  2613 => x"0cfe117e",
  2614 => x"29770580",
  2615 => x"eda00c52",
  2616 => x"59524354",
  2617 => x"5e515259",
  2618 => x"525d5759",
  2619 => x"5780d2c9",
  2620 => x"0480e792",
  2621 => x"0b80f52d",
  2622 => x"80e7910b",
  2623 => x"80f52d71",
  2624 => x"82802905",
  2625 => x"7080ed90",
  2626 => x"0c70a029",
  2627 => x"83ff0570",
  2628 => x"892a7080",
  2629 => x"eda40c80",
  2630 => x"e7970b80",
  2631 => x"f52d80e7",
  2632 => x"960b80f5",
  2633 => x"2d718280",
  2634 => x"29057080",
  2635 => x"edac0c7b",
  2636 => x"71291e70",
  2637 => x"80eda00c",
  2638 => x"7d80ed9c",
  2639 => x"0c730580",
  2640 => x"ed980c55",
  2641 => x"5e515155",
  2642 => x"55805180",
  2643 => x"cb8b2d81",
  2644 => x"557480e6",
  2645 => x"8c0c02a8",
  2646 => x"050d0402",
  2647 => x"ec050d76",
  2648 => x"70872c71",
  2649 => x"80ff0655",
  2650 => x"565480ed",
  2651 => x"8c088a38",
  2652 => x"73882c74",
  2653 => x"81ff0654",
  2654 => x"5580e780",
  2655 => x"5280ed94",
  2656 => x"08155180",
  2657 => x"c9a22d80",
  2658 => x"e68c0854",
  2659 => x"80e68c08",
  2660 => x"802ebb38",
  2661 => x"80ed8c08",
  2662 => x"802e9c38",
  2663 => x"72842980",
  2664 => x"e7800570",
  2665 => x"08525380",
  2666 => x"d9952d80",
  2667 => x"e68c08f0",
  2668 => x"0a065380",
  2669 => x"d3cc0472",
  2670 => x"1080e780",
  2671 => x"057080e0",
  2672 => x"2d525380",
  2673 => x"d9c62d80",
  2674 => x"e68c0853",
  2675 => x"72547380",
  2676 => x"e68c0c02",
  2677 => x"94050d04",
  2678 => x"02e0050d",
  2679 => x"7970842c",
  2680 => x"80edb408",
  2681 => x"05718f06",
  2682 => x"52555372",
  2683 => x"8b3880e7",
  2684 => x"80527351",
  2685 => x"80c9a22d",
  2686 => x"72a02980",
  2687 => x"e7800554",
  2688 => x"807480f5",
  2689 => x"2d565374",
  2690 => x"732e8338",
  2691 => x"81537481",
  2692 => x"e52e81f5",
  2693 => x"38817074",
  2694 => x"06545872",
  2695 => x"802e81e9",
  2696 => x"388b1480",
  2697 => x"f52d7083",
  2698 => x"2a790658",
  2699 => x"56769c38",
  2700 => x"80e4d008",
  2701 => x"53728938",
  2702 => x"7280eb80",
  2703 => x"0b81b72d",
  2704 => x"7680e4d0",
  2705 => x"0c735380",
  2706 => x"d68b0475",
  2707 => x"8f2e0981",
  2708 => x"0681b638",
  2709 => x"749f068d",
  2710 => x"2980eaf3",
  2711 => x"11515381",
  2712 => x"1480f52d",
  2713 => x"73708105",
  2714 => x"5581b72d",
  2715 => x"831480f5",
  2716 => x"2d737081",
  2717 => x"055581b7",
  2718 => x"2d851480",
  2719 => x"f52d7370",
  2720 => x"81055581",
  2721 => x"b72d8714",
  2722 => x"80f52d73",
  2723 => x"70810555",
  2724 => x"81b72d89",
  2725 => x"1480f52d",
  2726 => x"73708105",
  2727 => x"5581b72d",
  2728 => x"8e1480f5",
  2729 => x"2d737081",
  2730 => x"055581b7",
  2731 => x"2d901480",
  2732 => x"f52d7370",
  2733 => x"81055581",
  2734 => x"b72d9214",
  2735 => x"80f52d73",
  2736 => x"70810555",
  2737 => x"81b72d94",
  2738 => x"1480f52d",
  2739 => x"73708105",
  2740 => x"5581b72d",
  2741 => x"961480f5",
  2742 => x"2d737081",
  2743 => x"055581b7",
  2744 => x"2d981480",
  2745 => x"f52d7370",
  2746 => x"81055581",
  2747 => x"b72d9c14",
  2748 => x"80f52d73",
  2749 => x"70810555",
  2750 => x"81b72d9e",
  2751 => x"1480f52d",
  2752 => x"7381b72d",
  2753 => x"7780e4d0",
  2754 => x"0c805372",
  2755 => x"80e68c0c",
  2756 => x"02a0050d",
  2757 => x"0402cc05",
  2758 => x"0d7e605e",
  2759 => x"5a800b80",
  2760 => x"edb00880",
  2761 => x"edb40859",
  2762 => x"5c568058",
  2763 => x"80ed9008",
  2764 => x"782e81be",
  2765 => x"38778f06",
  2766 => x"a0175754",
  2767 => x"73923880",
  2768 => x"e7805276",
  2769 => x"51811757",
  2770 => x"80c9a22d",
  2771 => x"80e78056",
  2772 => x"807680f5",
  2773 => x"2d565474",
  2774 => x"742e8338",
  2775 => x"81547481",
  2776 => x"e52e8182",
  2777 => x"38817075",
  2778 => x"06555c73",
  2779 => x"802e80f6",
  2780 => x"388b1680",
  2781 => x"f52d9806",
  2782 => x"597880ea",
  2783 => x"388b537c",
  2784 => x"52755180",
  2785 => x"caca2d80",
  2786 => x"e68c0880",
  2787 => x"d9389c16",
  2788 => x"085180d9",
  2789 => x"952d80e6",
  2790 => x"8c08841b",
  2791 => x"0c9a1680",
  2792 => x"e02d5180",
  2793 => x"d9c62d80",
  2794 => x"e68c0880",
  2795 => x"e68c0888",
  2796 => x"1c0c80e6",
  2797 => x"8c085555",
  2798 => x"80ed8c08",
  2799 => x"802e9a38",
  2800 => x"941680e0",
  2801 => x"2d5180d9",
  2802 => x"c62d80e6",
  2803 => x"8c08902b",
  2804 => x"83fff00a",
  2805 => x"06701651",
  2806 => x"5473881b",
  2807 => x"0c787a0c",
  2808 => x"7b5480d8",
  2809 => x"b0048118",
  2810 => x"5880ed90",
  2811 => x"087826fe",
  2812 => x"c43880ed",
  2813 => x"8c08802e",
  2814 => x"b5387a51",
  2815 => x"80d2db2d",
  2816 => x"80e68c08",
  2817 => x"80e68c08",
  2818 => x"80ffffff",
  2819 => x"f806555b",
  2820 => x"7380ffff",
  2821 => x"fff82e96",
  2822 => x"3880e68c",
  2823 => x"08fe0580",
  2824 => x"ed840829",
  2825 => x"80ed9808",
  2826 => x"055780d6",
  2827 => x"aa048054",
  2828 => x"7380e68c",
  2829 => x"0c02b405",
  2830 => x"0d0402f4",
  2831 => x"050d7470",
  2832 => x"08810571",
  2833 => x"0c700880",
  2834 => x"ed880806",
  2835 => x"53537190",
  2836 => x"38881308",
  2837 => x"5180d2db",
  2838 => x"2d80e68c",
  2839 => x"0888140c",
  2840 => x"810b80e6",
  2841 => x"8c0c028c",
  2842 => x"050d0402",
  2843 => x"f0050d75",
  2844 => x"881108fe",
  2845 => x"0580ed84",
  2846 => x"082980ed",
  2847 => x"98081172",
  2848 => x"0880ed88",
  2849 => x"08060579",
  2850 => x"55535454",
  2851 => x"80c9a22d",
  2852 => x"0290050d",
  2853 => x"0402f405",
  2854 => x"0d747088",
  2855 => x"2a83fe80",
  2856 => x"06707298",
  2857 => x"2a077288",
  2858 => x"2b87fc80",
  2859 => x"80067398",
  2860 => x"2b81f00a",
  2861 => x"06717307",
  2862 => x"0780e68c",
  2863 => x"0c565153",
  2864 => x"51028c05",
  2865 => x"0d0402f8",
  2866 => x"050d028e",
  2867 => x"0580f52d",
  2868 => x"74882b07",
  2869 => x"7083ffff",
  2870 => x"0680e68c",
  2871 => x"0c510288",
  2872 => x"050d0402",
  2873 => x"f4050d74",
  2874 => x"76785354",
  2875 => x"52807125",
  2876 => x"97387270",
  2877 => x"81055480",
  2878 => x"f52d7270",
  2879 => x"81055481",
  2880 => x"b72dff11",
  2881 => x"5170eb38",
  2882 => x"807281b7",
  2883 => x"2d028c05",
  2884 => x"0d0402e8",
  2885 => x"050d7756",
  2886 => x"80705654",
  2887 => x"737624b7",
  2888 => x"3880ed90",
  2889 => x"08742eaf",
  2890 => x"38735180",
  2891 => x"d3d82d80",
  2892 => x"e68c0880",
  2893 => x"e68c0809",
  2894 => x"81057080",
  2895 => x"e68c0807",
  2896 => x"9f2a7705",
  2897 => x"81175757",
  2898 => x"53537476",
  2899 => x"24893880",
  2900 => x"ed900874",
  2901 => x"26d33872",
  2902 => x"80e68c0c",
  2903 => x"0298050d",
  2904 => x"0402f005",
  2905 => x"0d80e688",
  2906 => x"08165180",
  2907 => x"da922d80",
  2908 => x"e68c0880",
  2909 => x"2ea0388b",
  2910 => x"5380e68c",
  2911 => x"085280eb",
  2912 => x"805180d9",
  2913 => x"e32d80ed",
  2914 => x"bc085473",
  2915 => x"802e8738",
  2916 => x"80eb8051",
  2917 => x"732d0290",
  2918 => x"050d0402",
  2919 => x"dc050d80",
  2920 => x"705a5574",
  2921 => x"80e68808",
  2922 => x"25b53880",
  2923 => x"ed900875",
  2924 => x"2ead3878",
  2925 => x"5180d3d8",
  2926 => x"2d80e68c",
  2927 => x"08098105",
  2928 => x"7080e68c",
  2929 => x"08079f2a",
  2930 => x"7605811b",
  2931 => x"5b565474",
  2932 => x"80e68808",
  2933 => x"25893880",
  2934 => x"ed900879",
  2935 => x"26d53880",
  2936 => x"557880ed",
  2937 => x"90082781",
  2938 => x"e4387851",
  2939 => x"80d3d82d",
  2940 => x"80e68c08",
  2941 => x"802e81b4",
  2942 => x"3880e68c",
  2943 => x"088b0580",
  2944 => x"f52d7084",
  2945 => x"2a708106",
  2946 => x"77107884",
  2947 => x"2b80eb80",
  2948 => x"0b80f52d",
  2949 => x"5c5c5351",
  2950 => x"55567380",
  2951 => x"2e80ce38",
  2952 => x"7416822b",
  2953 => x"80ddf10b",
  2954 => x"80e4dc12",
  2955 => x"0c547775",
  2956 => x"311080ed",
  2957 => x"c0115556",
  2958 => x"90747081",
  2959 => x"055681b7",
  2960 => x"2da07481",
  2961 => x"b72d7681",
  2962 => x"ff068116",
  2963 => x"58547380",
  2964 => x"2e8b389c",
  2965 => x"5380eb80",
  2966 => x"5280dce4",
  2967 => x"048b5380",
  2968 => x"e68c0852",
  2969 => x"80edc216",
  2970 => x"5180dda2",
  2971 => x"04741682",
  2972 => x"2b80dae1",
  2973 => x"0b80e4dc",
  2974 => x"120c5476",
  2975 => x"81ff0681",
  2976 => x"16585473",
  2977 => x"802e8b38",
  2978 => x"9c5380eb",
  2979 => x"805280dd",
  2980 => x"99048b53",
  2981 => x"80e68c08",
  2982 => x"52777531",
  2983 => x"1080edc0",
  2984 => x"05517655",
  2985 => x"80d9e32d",
  2986 => x"80ddc104",
  2987 => x"74902975",
  2988 => x"31701080",
  2989 => x"edc00551",
  2990 => x"5480e68c",
  2991 => x"087481b7",
  2992 => x"2d811959",
  2993 => x"748b24a4",
  2994 => x"3880dbe1",
  2995 => x"04749029",
  2996 => x"75317010",
  2997 => x"80edc005",
  2998 => x"8c773157",
  2999 => x"51548074",
  3000 => x"81b72d9e",
  3001 => x"14ff1656",
  3002 => x"5474f338",
  3003 => x"02a4050d",
  3004 => x"0402fc05",
  3005 => x"0d80e688",
  3006 => x"08135180",
  3007 => x"da922d80",
  3008 => x"e68c0880",
  3009 => x"2e8a3880",
  3010 => x"e68c0851",
  3011 => x"80cb8b2d",
  3012 => x"800b80e6",
  3013 => x"880c80db",
  3014 => x"9b2db7e5",
  3015 => x"2d028405",
  3016 => x"0d0402fc",
  3017 => x"050d7251",
  3018 => x"70fd2eb2",
  3019 => x"3870fd24",
  3020 => x"8b3870fc",
  3021 => x"2e80d038",
  3022 => x"80df9104",
  3023 => x"70fe2eb9",
  3024 => x"3870ff2e",
  3025 => x"09810680",
  3026 => x"c83880e6",
  3027 => x"88085170",
  3028 => x"802ebe38",
  3029 => x"ff1180e6",
  3030 => x"880c80df",
  3031 => x"910480e6",
  3032 => x"8808f005",
  3033 => x"7080e688",
  3034 => x"0c517080",
  3035 => x"25a33880",
  3036 => x"0b80e688",
  3037 => x"0c80df91",
  3038 => x"0480e688",
  3039 => x"08810580",
  3040 => x"e6880c80",
  3041 => x"df910480",
  3042 => x"e6880890",
  3043 => x"0580e688",
  3044 => x"0c80db9b",
  3045 => x"2db7e52d",
  3046 => x"0284050d",
  3047 => x"0402fc05",
  3048 => x"0d800b80",
  3049 => x"e6880c80",
  3050 => x"db9b2db6",
  3051 => x"ee2d80e6",
  3052 => x"8c0880e5",
  3053 => x"f80c80e4",
  3054 => x"d451b98b",
  3055 => x"2d028405",
  3056 => x"0d047180",
  3057 => x"edbc0c04",
  3058 => x"00ffffff",
  3059 => x"ff00ffff",
  3060 => x"ffff00ff",
  3061 => x"ffffff00",
  3062 => x"52657365",
  3063 => x"74205369",
  3064 => x"6e636c61",
  3065 => x"69722051",
  3066 => x"4c000000",
  3067 => x"5363616e",
  3068 => x"6c696e65",
  3069 => x"73000000",
  3070 => x"4d6f756e",
  3071 => x"74204d44",
  3072 => x"56201000",
  3073 => x"45786974",
  3074 => x"00000000",
  3075 => x"56696465",
  3076 => x"6f205041",
  3077 => x"4c200000",
  3078 => x"56696465",
  3079 => x"6f204e54",
  3080 => x"53430000",
  3081 => x"52414d20",
  3082 => x"3132386b",
  3083 => x"62000000",
  3084 => x"52414d20",
  3085 => x"3634306b",
  3086 => x"62000000",
  3087 => x"4d445620",
  3088 => x"6e6f726d",
  3089 => x"616c2020",
  3090 => x"00000000",
  3091 => x"4d445620",
  3092 => x"72657665",
  3093 => x"72736564",
  3094 => x"00000000",
  3095 => x"524f4d20",
  3096 => x"6c6f6164",
  3097 => x"696e6720",
  3098 => x"6661696c",
  3099 => x"65640000",
  3100 => x"4f4b0000",
  3101 => x"496e6974",
  3102 => x"69616c69",
  3103 => x"7a696e67",
  3104 => x"20534420",
  3105 => x"63617264",
  3106 => x"0a000000",
  3107 => x"4c6f6164",
  3108 => x"696e6720",
  3109 => x"514c2e52",
  3110 => x"4f4d2e2e",
  3111 => x"2e0a0000",
  3112 => x"514c2020",
  3113 => x"20202020",
  3114 => x"524f4d00",
  3115 => x"16200000",
  3116 => x"14200000",
  3117 => x"15200000",
  3118 => x"53442069",
  3119 => x"6e69742e",
  3120 => x"2e2e0a00",
  3121 => x"53442063",
  3122 => x"61726420",
  3123 => x"72657365",
  3124 => x"74206661",
  3125 => x"696c6564",
  3126 => x"210a0000",
  3127 => x"53444843",
  3128 => x"20657272",
  3129 => x"6f72210a",
  3130 => x"00000000",
  3131 => x"57726974",
  3132 => x"65206661",
  3133 => x"696c6564",
  3134 => x"0a000000",
  3135 => x"52656164",
  3136 => x"20666169",
  3137 => x"6c65640a",
  3138 => x"00000000",
  3139 => x"43617264",
  3140 => x"20696e69",
  3141 => x"74206661",
  3142 => x"696c6564",
  3143 => x"0a000000",
  3144 => x"46415431",
  3145 => x"36202020",
  3146 => x"00000000",
  3147 => x"46415433",
  3148 => x"32202020",
  3149 => x"00000000",
  3150 => x"4e6f2070",
  3151 => x"61727469",
  3152 => x"74696f6e",
  3153 => x"20736967",
  3154 => x"0a000000",
  3155 => x"42616420",
  3156 => x"70617274",
  3157 => x"0a000000",
  3158 => x"4261636b",
  3159 => x"00000000",
  3160 => x"00000002",
  3161 => x"00000002",
  3162 => x"00002fd8",
  3163 => x"0000035a",
  3164 => x"00000003",
  3165 => x"000031d4",
  3166 => x"00000002",
  3167 => x"00000003",
  3168 => x"000031cc",
  3169 => x"00000002",
  3170 => x"00000003",
  3171 => x"000031c4",
  3172 => x"00000002",
  3173 => x"00000001",
  3174 => x"00002fec",
  3175 => x"00000005",
  3176 => x"00000002",
  3177 => x"00002ff8",
  3178 => x"00002f9d",
  3179 => x"00000002",
  3180 => x"00003004",
  3181 => x"00001b8b",
  3182 => x"00000000",
  3183 => x"00000000",
  3184 => x"00000000",
  3185 => x"0000300c",
  3186 => x"00003018",
  3187 => x"00003024",
  3188 => x"00003030",
  3189 => x"0000303c",
  3190 => x"0000304c",
  3191 => x"00000004",
  3192 => x"0000305c",
  3193 => x"000031dc",
  3194 => x"00000004",
  3195 => x"00003070",
  3196 => x"00003164",
  3197 => x"00000000",
  3198 => x"00000000",
  3199 => x"00000000",
  3200 => x"00000000",
  3201 => x"00000000",
  3202 => x"00000000",
  3203 => x"00000000",
  3204 => x"00000000",
  3205 => x"00000000",
  3206 => x"00000000",
  3207 => x"00000000",
  3208 => x"00000000",
  3209 => x"00000000",
  3210 => x"00000000",
  3211 => x"00000000",
  3212 => x"00000000",
  3213 => x"00000000",
  3214 => x"00000000",
  3215 => x"00000000",
  3216 => x"00000000",
  3217 => x"00000000",
  3218 => x"00000000",
  3219 => x"00000000",
  3220 => x"00000000",
  3221 => x"00000002",
  3222 => x"000036c0",
  3223 => x"00002d61",
  3224 => x"00000002",
  3225 => x"000036de",
  3226 => x"00002d61",
  3227 => x"00000002",
  3228 => x"000036fc",
  3229 => x"00002d61",
  3230 => x"00000002",
  3231 => x"0000371a",
  3232 => x"00002d61",
  3233 => x"00000002",
  3234 => x"00003738",
  3235 => x"00002d61",
  3236 => x"00000002",
  3237 => x"00003756",
  3238 => x"00002d61",
  3239 => x"00000002",
  3240 => x"00003774",
  3241 => x"00002d61",
  3242 => x"00000002",
  3243 => x"00003792",
  3244 => x"00002d61",
  3245 => x"00000002",
  3246 => x"000037b0",
  3247 => x"00002d61",
  3248 => x"00000002",
  3249 => x"000037ce",
  3250 => x"00002d61",
  3251 => x"00000002",
  3252 => x"000037ec",
  3253 => x"00002d61",
  3254 => x"00000002",
  3255 => x"0000380a",
  3256 => x"00002d61",
  3257 => x"00000002",
  3258 => x"00003828",
  3259 => x"00002d61",
  3260 => x"00000004",
  3261 => x"00003158",
  3262 => x"00000000",
  3263 => x"00000000",
  3264 => x"00000000",
  3265 => x"00002f22",
  3266 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

