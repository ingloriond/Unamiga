library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom_t49 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(10 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom_t49 is
	type rom is array(0 to  2047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"04",X"09",X"00",X"04",X"DE",X"00",X"00",X"24",X"00",X"65",X"15",X"35",X"85",X"95",X"8A",X"01",
		X"9A",X"FD",X"8A",X"04",X"8A",X"08",X"8A",X"10",X"8A",X"20",X"8A",X"40",X"8A",X"80",X"B8",X"20",
		X"BA",X"60",X"B0",X"00",X"18",X"EA",X"22",X"B8",X"29",X"B0",X"FF",X"B8",X"2B",X"B0",X"2C",X"B8",
		X"24",X"B0",X"03",X"B8",X"4E",X"B0",X"52",X"18",X"B0",X"52",X"18",X"B0",X"69",X"18",X"B0",X"69",
		X"A5",X"14",X"4A",X"0A",X"53",X"80",X"C6",X"43",X"A4",X"00",X"65",X"D5",X"B8",X"20",X"F0",X"53",
		X"02",X"B8",X"22",X"C6",X"5D",X"F0",X"43",X"04",X"53",X"EF",X"A0",X"64",X"E4",X"BA",X"00",X"B8",
		X"4C",X"F0",X"37",X"17",X"53",X"3F",X"03",X"EC",X"E6",X"6E",X"FA",X"43",X"10",X"AA",X"18",X"F0",
		X"37",X"17",X"53",X"3F",X"03",X"EC",X"E6",X"7C",X"FA",X"43",X"20",X"AA",X"FA",X"37",X"B8",X"20",
		X"50",X"B8",X"22",X"92",X"9F",X"B2",X"91",X"65",X"23",X"00",X"62",X"35",X"25",X"55",X"FF",X"C5",
		X"93",X"F0",X"43",X"01",X"A0",X"BA",X"51",X"B9",X"4D",X"BE",X"80",X"BC",X"80",X"04",X"B4",X"B2",
		X"AF",X"F0",X"53",X"FE",X"A0",X"BA",X"4F",X"B9",X"4C",X"BE",X"97",X"BC",X"40",X"04",X"B4",X"F0",
		X"12",X"A1",X"04",X"91",X"FC",X"37",X"50",X"53",X"FD",X"43",X"08",X"A0",X"C8",X"B0",X"00",X"18",
		X"18",X"B0",X"00",X"B8",X"4B",X"FA",X"A0",X"A8",X"F0",X"AA",X"B8",X"22",X"B5",X"BB",X"00",X"05",
		X"35",X"FC",X"F2",X"D9",X"FF",X"C5",X"9A",X"EF",X"93",X"FF",X"C5",X"9A",X"DF",X"93",X"B6",X"E1",
		X"93",X"D5",X"AF",X"23",X"FF",X"62",X"25",X"45",X"15",X"FF",X"93",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B6",X"03",X"93",X"D5",X"AF",X"65",X"23",X"FC",X"62",X"45",X"76",X"37",X"B8",X"22",X"F0",X"53",
		X"04",X"96",X"15",X"04",X"4A",X"64",X"27",X"B8",X"20",X"12",X"21",X"F0",X"43",X"10",X"A0",X"A4",
		X"00",X"F0",X"43",X"20",X"A0",X"A4",X"00",X"B8",X"20",X"12",X"31",X"F0",X"53",X"EF",X"A0",X"A4",
		X"00",X"F0",X"53",X"DF",X"A0",X"A4",X"00",X"0A",X"53",X"01",X"2B",X"96",X"55",X"2B",X"96",X"4C",
		X"F0",X"53",X"F7",X"A0",X"C8",X"B0",X"00",X"18",X"BB",X"09",X"FF",X"93",X"65",X"35",X"05",X"F0",
		X"43",X"08",X"A0",X"FF",X"93",X"2B",X"EB",X"8A",X"65",X"35",X"05",X"96",X"64",X"F0",X"5C",X"96",
		X"84",X"FC",X"40",X"A0",X"FA",X"A8",X"FD",X"A0",X"F1",X"07",X"A1",X"18",X"F8",X"6E",X"F8",X"E6",
		X"73",X"03",X"E9",X"AA",X"B8",X"22",X"F1",X"03",X"14",X"96",X"81",X"8A",X"30",X"F0",X"43",X"02",
		X"A0",X"18",X"10",X"C8",X"F0",X"43",X"08",X"A0",X"FF",X"93",X"67",X"FD",X"67",X"AD",X"FF",X"93",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"53",X"80",X"C6",X"07",X"A4",X"00",X"F4",X"4F",X"03",X"0C",X"B3",X"1C",X"28",X"1E",X"1E",
		X"20",X"20",X"89",X"89",X"4D",X"76",X"22",X"24",X"C3",X"CF",X"E3",X"F0",X"04",X"09",X"24",X"17",
		X"24",X"27",X"64",X"00",X"64",X"1F",X"A4",X"00",X"0A",X"53",X"40",X"B8",X"20",X"40",X"53",X"CF",
		X"72",X"34",X"44",X"36",X"43",X"01",X"AA",X"B8",X"4C",X"F0",X"C6",X"40",X"FA",X"43",X"10",X"AA",
		X"18",X"F0",X"C6",X"48",X"FA",X"43",X"20",X"AA",X"FA",X"F4",X"84",X"A4",X"00",X"B8",X"2B",X"F0",
		X"03",X"D4",X"97",X"67",X"AA",X"B9",X"20",X"F1",X"53",X"08",X"4A",X"F4",X"89",X"FA",X"C6",X"6E",
		X"B9",X"2C",X"F1",X"F4",X"89",X"19",X"F1",X"F4",X"84",X"19",X"EA",X"62",X"B0",X"2C",X"B8",X"20",
		X"F0",X"53",X"FE",X"A0",X"A4",X"00",X"F4",X"4F",X"53",X"07",X"17",X"AA",X"23",X"00",X"97",X"A7",
		X"F7",X"EA",X"80",X"B4",X"C8",X"F4",X"84",X"A4",X"00",X"12",X"93",X"B8",X"4C",X"BC",X"97",X"BD",
		X"4E",X"44",X"99",X"B8",X"4D",X"BC",X"80",X"BD",X"50",X"F0",X"37",X"17",X"53",X"3F",X"AB",X"B9",
		X"22",X"F1",X"53",X"C0",X"4B",X"F4",X"84",X"FB",X"C6",X"C1",X"FD",X"A9",X"F1",X"A9",X"F1",X"F4",
		X"84",X"10",X"19",X"F9",X"6C",X"E6",X"BB",X"F9",X"03",X"E9",X"A9",X"EB",X"AE",X"FD",X"A8",X"F9",
		X"A0",X"A4",X"00",X"F4",X"4F",X"12",X"CB",X"9A",X"F7",X"A4",X"00",X"8A",X"08",X"A4",X"00",X"F4",
		X"4F",X"53",X"07",X"03",X"DB",X"A3",X"B8",X"24",X"A0",X"A4",X"00",X"01",X"03",X"07",X"0F",X"1F",
		X"3F",X"7F",X"FF",X"F4",X"3A",X"B9",X"25",X"F1",X"F4",X"84",X"19",X"F1",X"F4",X"84",X"A4",X"00",
		X"F4",X"7C",X"F4",X"84",X"A4",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B8",X"3A",X"B9",X"08",X"F4",X"7C",X"A0",X"18",X"E9",X"04",X"94",X"15",X"18",X"A0",X"18",X"A0",
		X"B9",X"05",X"18",X"B0",X"00",X"E9",X"12",X"B8",X"20",X"F0",X"43",X"02",X"A0",X"A4",X"00",X"B8",
		X"20",X"F0",X"53",X"FD",X"A0",X"A4",X"00",X"65",X"B8",X"20",X"F0",X"53",X"02",X"96",X"3B",X"B8",
		X"22",X"F0",X"53",X"FB",X"53",X"DF",X"A0",X"9A",X"FD",X"04",X"4A",X"B8",X"3E",X"F0",X"96",X"44",
		X"18",X"F0",X"C6",X"65",X"B8",X"4A",X"10",X"10",X"B9",X"47",X"B8",X"44",X"F0",X"96",X"51",X"23",
		X"FF",X"F4",X"16",X"B8",X"4A",X"F0",X"F4",X"16",X"B8",X"3F",X"19",X"F4",X"0B",X"E6",X"65",X"B8",
		X"22",X"F0",X"43",X"20",X"A0",X"B9",X"45",X"B8",X"44",X"F0",X"96",X"6E",X"23",X"FF",X"F4",X"16",
		X"B8",X"4A",X"F0",X"F4",X"16",X"B8",X"3D",X"19",X"F4",X"0B",X"E6",X"E4",X"B8",X"4A",X"F0",X"03",
		X"03",X"A0",X"B8",X"45",X"B0",X"00",X"18",X"B0",X"00",X"B8",X"42",X"B9",X"40",X"F1",X"47",X"43",
		X"F0",X"72",X"95",X"53",X"0F",X"60",X"A0",X"B9",X"3A",X"F4",X"00",X"F6",X"A5",X"B9",X"3B",X"F4",
		X"00",X"C6",X"A5",X"F6",X"D3",X"B8",X"4A",X"10",X"10",X"B8",X"40",X"F0",X"B8",X"49",X"43",X"F0",
		X"17",X"C6",X"BD",X"07",X"53",X"0F",X"C6",X"C2",X"37",X"17",X"60",X"F6",X"C2",X"10",X"94",X"15",
		X"64",X"D3",X"B0",X"00",X"B9",X"40",X"F1",X"47",X"37",X"17",X"53",X"0F",X"47",X"AA",X"F1",X"53",
		X"0F",X"4A",X"A1",X"B9",X"41",X"F1",X"47",X"A1",X"94",X"22",X"B9",X"42",X"61",X"19",X"A1",X"B9",
		X"41",X"F1",X"47",X"A1",X"B8",X"22",X"F0",X"53",X"10",X"C6",X"F3",X"9A",X"FD",X"F0",X"53",X"EF",
		X"A0",X"84",X"00",X"8A",X"02",X"F0",X"43",X"10",X"A0",X"84",X"00",X"00",X"00",X"00",X"00",X"00",
		X"94",X"22",X"B9",X"43",X"61",X"19",X"A1",X"37",X"17",X"65",X"62",X"35",X"25",X"55",X"B8",X"4A",
		X"B0",X"04",X"FF",X"C5",X"93",X"B8",X"40",X"F0",X"B9",X"3B",X"F2",X"1D",X"C9",X"B8",X"42",X"F1",
		X"A0",X"83",X"B8",X"41",X"F0",X"72",X"29",X"27",X"83",X"B8",X"4A",X"F0",X"03",X"07",X"A0",X"F4",
		X"3A",X"B8",X"41",X"B9",X"25",X"F0",X"53",X"07",X"17",X"AA",X"27",X"97",X"A7",X"F7",X"EA",X"3C",
		X"51",X"83",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"B8",X"27",X"10",X"BA",X"08",X"23",X"80",X"B4",X"C8",X"AE",X"53",X"07",X"03",X"C0",X"A3",X"AC",
		X"B8",X"28",X"D0",X"C6",X"21",X"B9",X"20",X"F1",X"43",X"04",X"53",X"F7",X"A1",X"FC",X"A0",X"A4",
		X"BE",X"FE",X"53",X"F8",X"BE",X"FF",X"B4",X"D3",X"F6",X"3F",X"CA",X"FB",X"77",X"B4",X"C8",X"B4",
		X"D3",X"F6",X"3F",X"EA",X"2B",X"FE",X"17",X"96",X"4E",X"B8",X"20",X"F0",X"53",X"FB",X"A0",X"B8",
		X"20",X"F0",X"53",X"F7",X"A0",X"B8",X"29",X"B0",X"FF",X"18",X"B0",X"00",X"A4",X"BE",X"B8",X"20",
		X"F0",X"53",X"04",X"96",X"BE",X"B8",X"29",X"F0",X"DE",X"C6",X"62",X"FE",X"A0",X"18",X"B0",X"00",
		X"A4",X"BE",X"18",X"F0",X"03",X"FC",X"C6",X"6D",X"F6",X"B8",X"10",X"A4",X"BE",X"10",X"B8",X"28",
		X"F0",X"03",X"FD",X"96",X"8D",X"FE",X"03",X"C1",X"96",X"8D",X"9A",X"FB",X"15",X"35",X"65",X"8A",
		X"10",X"8A",X"20",X"B8",X"FF",X"B9",X"FF",X"E9",X"87",X"E8",X"85",X"04",X"09",X"B8",X"2B",X"F0",
		X"A9",X"03",X"C6",X"C6",X"B0",X"B8",X"28",X"F0",X"A1",X"19",X"FE",X"A1",X"19",X"F9",X"B8",X"2B",
		X"A0",X"B8",X"20",X"F0",X"43",X"01",X"A0",X"B8",X"27",X"F0",X"B9",X"25",X"F4",X"16",X"A4",X"BE",
		X"B8",X"38",X"F0",X"43",X"08",X"A0",X"A4",X"BE",X"B8",X"20",X"F0",X"43",X"08",X"A0",X"C4",X"00",
		X"00",X"04",X"02",X"06",X"01",X"05",X"03",X"07",X"39",X"AB",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"08",X"93",X"C6",X"F9",X"2E",X"17",X"C6",X"DC",X"97",X"A7",X"83",X"BC",X"08",X"FE",X"F2",
		X"E8",X"E7",X"EC",X"DF",X"BE",X"FF",X"97",X"83",X"53",X"7F",X"96",X"D9",X"FA",X"07",X"37",X"53",
		X"07",X"E7",X"E7",X"E7",X"AE",X"FC",X"07",X"4E",X"AE",X"97",X"83",X"00",X"00",X"00",X"00",X"00",
		X"76",X"11",X"B8",X"22",X"F0",X"53",X"20",X"C6",X"0F",X"B8",X"20",X"F0",X"53",X"FD",X"A0",X"44",
		X"00",X"B8",X"22",X"F0",X"53",X"08",X"C6",X"4A",X"B8",X"24",X"B9",X"21",X"11",X"F4",X"00",X"E6",
		X"4A",X"B8",X"20",X"F0",X"53",X"80",X"C6",X"3E",X"85",X"F0",X"53",X"7F",X"A0",X"65",X"15",X"35",
		X"B5",X"D5",X"B8",X"4B",X"F0",X"A9",X"FA",X"A1",X"C5",X"14",X"4A",X"95",X"44",X"00",X"8A",X"30",
		X"B8",X"20",X"F0",X"43",X"80",X"A0",X"B1",X"00",X"44",X"00",X"B9",X"23",X"F1",X"03",X"E9",X"F6",
		X"3E",X"B8",X"22",X"F0",X"53",X"02",X"96",X"3E",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"C6",X"07",X"37",X"17",X"61",X"83",X"F1",X"97",X"A7",X"83",X"F4",X"00",X"96",X"15",X"C8",
		X"C9",X"F4",X"00",X"18",X"19",X"83",X"61",X"A1",X"19",X"23",X"00",X"71",X"A1",X"C9",X"83",X"BD",
		X"00",X"BE",X"00",X"97",X"B8",X"08",X"FA",X"67",X"AA",X"E6",X"31",X"FB",X"6D",X"AD",X"FC",X"7E",
		X"AE",X"FB",X"F7",X"AB",X"FC",X"F7",X"AC",X"E8",X"26",X"83",X"B9",X"26",X"F1",X"AA",X"BB",X"8D",
		X"F4",X"1F",X"FE",X"B9",X"26",X"A1",X"C9",X"FD",X"F4",X"16",X"23",X"8B",X"F4",X"16",X"83",X"BE",
		X"00",X"BF",X"04",X"0A",X"53",X"80",X"96",X"53",X"90",X"0A",X"90",X"F7",X"FE",X"F7",X"AE",X"EF",
		X"53",X"93",X"BF",X"04",X"AE",X"0A",X"53",X"80",X"96",X"65",X"FE",X"90",X"F2",X"72",X"9A",X"7F",
		X"E4",X"74",X"8A",X"80",X"90",X"E7",X"AE",X"8A",X"80",X"EF",X"65",X"93",X"F4",X"4F",X"47",X"AD",
		X"F4",X"4F",X"4D",X"93",X"F4",X"62",X"F4",X"62",X"93",X"47",X"F4",X"62",X"93",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
